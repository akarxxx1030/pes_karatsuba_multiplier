module spm (iX,
    iY,
    oO);
 input [63:0] iX;
 input [63:0] iY;
 output [127:0] oO;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire _17588_;
 wire _17589_;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire _17625_;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire _17629_;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire _17652_;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire _17698_;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire _17703_;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire _17724_;
 wire _17725_;
 wire _17726_;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire _17762_;
 wire _17763_;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire _17778_;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire _17978_;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire _17988_;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire _17994_;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire _17999_;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire _18109_;
 wire _18110_;
 wire _18111_;
 wire _18112_;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire _18117_;
 wire _18118_;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire _18124_;
 wire _18125_;
 wire _18126_;
 wire _18127_;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire _18131_;
 wire _18132_;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire _18145_;
 wire _18146_;
 wire _18147_;
 wire _18148_;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire _18176_;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire _18180_;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire _18244_;
 wire _18245_;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire _18322_;
 wire _18323_;
 wire _18324_;
 wire _18325_;
 wire _18326_;
 wire _18327_;
 wire _18328_;
 wire _18329_;
 wire _18330_;
 wire _18331_;
 wire _18332_;
 wire _18333_;
 wire _18334_;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire _18338_;
 wire _18339_;
 wire _18340_;
 wire _18341_;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire _18354_;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire _18358_;
 wire _18359_;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire _18364_;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire _18368_;
 wire _18369_;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire _18378_;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire _18389_;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire _18396_;
 wire _18397_;
 wire _18398_;
 wire _18399_;
 wire _18400_;
 wire _18401_;
 wire _18402_;
 wire _18403_;
 wire _18404_;
 wire _18405_;
 wire _18406_;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire _18411_;
 wire _18412_;
 wire _18413_;
 wire _18414_;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire _18420_;
 wire _18421_;
 wire _18422_;
 wire _18423_;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire _18428_;
 wire _18429_;
 wire _18430_;
 wire _18431_;
 wire _18432_;
 wire _18433_;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire _18438_;
 wire _18439_;
 wire _18440_;
 wire _18441_;
 wire _18442_;
 wire _18443_;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire _18448_;
 wire _18449_;
 wire _18450_;
 wire _18451_;
 wire _18452_;
 wire _18453_;
 wire _18454_;
 wire _18455_;
 wire _18456_;
 wire _18457_;
 wire _18458_;
 wire _18459_;
 wire _18460_;
 wire _18461_;
 wire _18462_;
 wire _18463_;
 wire _18464_;
 wire _18465_;
 wire _18466_;
 wire _18467_;
 wire _18468_;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire _18472_;
 wire _18473_;
 wire _18474_;
 wire _18475_;
 wire _18476_;
 wire _18477_;
 wire _18478_;
 wire _18479_;
 wire _18480_;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire _18484_;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire _18491_;
 wire _18492_;
 wire _18493_;
 wire _18494_;
 wire _18495_;
 wire _18496_;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire _18504_;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire _18508_;
 wire _18509_;
 wire _18510_;
 wire _18511_;
 wire _18512_;
 wire _18513_;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire _18519_;
 wire _18520_;
 wire _18521_;
 wire _18522_;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire _18527_;
 wire _18528_;
 wire _18529_;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire _18534_;
 wire _18535_;
 wire _18536_;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire _18541_;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire _18546_;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire _18556_;
 wire _18557_;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire _18566_;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire _18580_;
 wire _18581_;
 wire _18582_;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire _18606_;
 wire _18607_;
 wire _18608_;
 wire _18609_;
 wire _18610_;
 wire _18611_;
 wire _18612_;
 wire _18613_;
 wire _18614_;
 wire _18615_;
 wire _18616_;
 wire _18617_;
 wire _18618_;
 wire _18619_;
 wire _18620_;
 wire _18621_;
 wire _18622_;
 wire _18623_;
 wire _18624_;
 wire _18625_;
 wire _18626_;
 wire _18627_;
 wire _18628_;
 wire _18629_;
 wire _18630_;
 wire _18631_;
 wire _18632_;
 wire _18633_;
 wire _18634_;
 wire _18635_;
 wire _18636_;
 wire _18637_;
 wire _18638_;
 wire _18639_;
 wire _18640_;
 wire _18641_;
 wire _18642_;
 wire _18643_;
 wire _18644_;
 wire _18645_;
 wire _18646_;
 wire _18647_;
 wire _18648_;
 wire _18649_;
 wire _18650_;
 wire _18651_;
 wire _18652_;
 wire _18653_;
 wire _18654_;
 wire _18655_;
 wire _18656_;
 wire _18657_;
 wire _18658_;
 wire _18659_;
 wire _18660_;
 wire _18661_;
 wire _18662_;
 wire _18663_;
 wire _18664_;
 wire _18665_;
 wire _18666_;
 wire _18667_;
 wire _18668_;
 wire _18669_;
 wire _18670_;
 wire _18671_;
 wire _18672_;
 wire _18673_;
 wire _18674_;
 wire _18675_;
 wire _18676_;
 wire _18677_;
 wire _18678_;
 wire _18679_;
 wire _18680_;
 wire _18681_;
 wire _18682_;
 wire _18683_;
 wire _18684_;
 wire _18685_;
 wire _18686_;
 wire _18687_;
 wire _18688_;
 wire _18689_;
 wire _18690_;
 wire _18691_;
 wire _18692_;
 wire _18693_;
 wire _18694_;
 wire _18695_;
 wire _18696_;
 wire _18697_;
 wire _18698_;
 wire _18699_;
 wire _18700_;
 wire _18701_;
 wire _18702_;
 wire _18703_;
 wire _18704_;
 wire _18705_;
 wire _18706_;
 wire _18707_;
 wire _18708_;
 wire _18709_;
 wire _18710_;
 wire _18711_;
 wire _18712_;
 wire _18713_;
 wire _18714_;
 wire _18715_;
 wire _18716_;
 wire _18717_;
 wire _18718_;
 wire _18719_;
 wire _18720_;
 wire _18721_;
 wire _18722_;
 wire _18723_;
 wire _18724_;
 wire _18725_;
 wire _18726_;
 wire _18727_;
 wire _18728_;
 wire _18729_;
 wire _18730_;
 wire _18731_;
 wire _18732_;
 wire _18733_;
 wire _18734_;
 wire _18735_;
 wire _18736_;
 wire _18737_;
 wire _18738_;
 wire _18739_;
 wire _18740_;
 wire _18741_;
 wire _18742_;
 wire _18743_;
 wire _18744_;
 wire _18745_;
 wire _18746_;
 wire _18747_;
 wire _18748_;
 wire _18749_;
 wire _18750_;
 wire _18751_;
 wire _18752_;
 wire _18753_;
 wire _18754_;
 wire _18755_;
 wire _18756_;
 wire _18757_;
 wire _18758_;
 wire _18759_;
 wire _18760_;
 wire _18761_;
 wire _18762_;
 wire _18763_;
 wire _18764_;
 wire _18765_;
 wire _18766_;
 wire _18767_;
 wire _18768_;
 wire _18769_;
 wire _18770_;
 wire _18771_;
 wire _18772_;
 wire _18773_;
 wire _18774_;
 wire _18775_;
 wire _18776_;
 wire _18777_;
 wire _18778_;
 wire _18779_;
 wire _18780_;
 wire _18781_;
 wire _18782_;
 wire _18783_;
 wire _18784_;
 wire _18785_;
 wire _18786_;
 wire _18787_;
 wire _18788_;
 wire _18789_;
 wire _18790_;
 wire _18791_;
 wire _18792_;
 wire _18793_;
 wire _18794_;
 wire _18795_;
 wire _18796_;
 wire _18797_;
 wire _18798_;
 wire _18799_;
 wire _18800_;
 wire _18801_;
 wire _18802_;
 wire _18803_;
 wire _18804_;
 wire _18805_;
 wire _18806_;
 wire _18807_;
 wire _18808_;
 wire _18809_;
 wire _18810_;
 wire _18811_;
 wire _18812_;
 wire _18813_;
 wire _18814_;
 wire _18815_;
 wire _18816_;
 wire _18817_;
 wire _18818_;
 wire _18819_;
 wire _18820_;
 wire _18821_;
 wire _18822_;
 wire _18823_;
 wire _18824_;
 wire _18825_;
 wire _18826_;
 wire _18827_;
 wire _18828_;
 wire _18829_;
 wire _18830_;
 wire _18831_;
 wire _18832_;
 wire _18833_;
 wire _18834_;
 wire _18835_;
 wire _18836_;
 wire _18837_;
 wire _18838_;
 wire _18839_;
 wire _18840_;
 wire _18841_;
 wire _18842_;
 wire _18843_;
 wire _18844_;
 wire _18845_;
 wire _18846_;
 wire _18847_;
 wire _18848_;
 wire _18849_;
 wire _18850_;
 wire _18851_;
 wire _18852_;
 wire _18853_;
 wire _18854_;
 wire _18855_;
 wire _18856_;
 wire _18857_;
 wire _18858_;
 wire _18859_;
 wire _18860_;
 wire _18861_;
 wire _18862_;
 wire _18863_;
 wire _18864_;
 wire _18865_;
 wire _18866_;
 wire _18867_;
 wire _18868_;
 wire _18869_;
 wire _18870_;
 wire _18871_;
 wire _18872_;
 wire _18873_;
 wire _18874_;
 wire _18875_;
 wire _18876_;
 wire _18877_;
 wire _18878_;
 wire _18879_;
 wire _18880_;
 wire _18881_;
 wire _18882_;
 wire _18883_;
 wire _18884_;
 wire _18885_;
 wire _18886_;
 wire _18887_;
 wire _18888_;
 wire _18889_;
 wire _18890_;
 wire _18891_;
 wire _18892_;
 wire _18893_;
 wire _18894_;
 wire _18895_;
 wire _18896_;
 wire _18897_;
 wire _18898_;
 wire _18899_;
 wire _18900_;
 wire _18901_;
 wire _18902_;
 wire _18903_;
 wire _18904_;
 wire _18905_;
 wire _18906_;
 wire _18907_;
 wire _18908_;
 wire _18909_;
 wire _18910_;
 wire _18911_;
 wire _18912_;
 wire _18913_;
 wire _18914_;
 wire _18915_;
 wire _18916_;
 wire _18917_;
 wire _18918_;
 wire _18919_;
 wire _18920_;
 wire _18921_;
 wire _18922_;
 wire _18923_;
 wire _18924_;
 wire _18925_;
 wire _18926_;
 wire _18927_;
 wire _18928_;
 wire _18929_;

 sky130_fd_sc_hd__nand2_2 _18930_ (.A(iY[0]),
    .B(iX[0]),
    .Y(_10801_));
 sky130_fd_sc_hd__inv_2 _18931_ (.A(_10801_),
    .Y(oO[0]));
 sky130_fd_sc_hd__a22oi_2 _18932_ (.A1(iY[0]),
    .A2(iX[1]),
    .B1(iY[1]),
    .B2(iX[0]),
    .Y(_10822_));
 sky130_fd_sc_hd__and3_2 _18933_ (.A(iX[1]),
    .B(iY[1]),
    .C(oO[0]),
    .X(_10832_));
 sky130_fd_sc_hd__or2_2 _18934_ (.A(_10822_),
    .B(_10832_),
    .X(_10843_));
 sky130_fd_sc_hd__inv_2 _18935_ (.A(_10843_),
    .Y(oO[1]));
 sky130_fd_sc_hd__and4_2 _18936_ (.A(iY[0]),
    .B(iX[1]),
    .C(iY[1]),
    .D(iX[2]),
    .X(_10864_));
 sky130_fd_sc_hd__a22oi_2 _18937_ (.A1(iX[1]),
    .A2(iY[1]),
    .B1(iX[2]),
    .B2(iY[0]),
    .Y(_10875_));
 sky130_fd_sc_hd__nor2_2 _18938_ (.A(_10864_),
    .B(_10875_),
    .Y(_10886_));
 sky130_fd_sc_hd__nand2_2 _18939_ (.A(iX[0]),
    .B(iY[2]),
    .Y(_10897_));
 sky130_fd_sc_hd__xnor2_2 _18940_ (.A(_10886_),
    .B(_10897_),
    .Y(_10908_));
 sky130_fd_sc_hd__nand2_2 _18941_ (.A(_10832_),
    .B(_10908_),
    .Y(_10919_));
 sky130_fd_sc_hd__or2_2 _18942_ (.A(_10832_),
    .B(_10908_),
    .X(_10930_));
 sky130_fd_sc_hd__and2_2 _18943_ (.A(_10919_),
    .B(_10930_),
    .X(_10941_));
 sky130_fd_sc_hd__buf_1 _18944_ (.A(_10941_),
    .X(oO[2]));
 sky130_fd_sc_hd__and4_2 _18945_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[2]),
    .D(iX[3]),
    .X(_10962_));
 sky130_fd_sc_hd__a22oi_2 _18946_ (.A1(iY[1]),
    .A2(iX[2]),
    .B1(iX[3]),
    .B2(iY[0]),
    .Y(_10973_));
 sky130_fd_sc_hd__nor2_2 _18947_ (.A(_10962_),
    .B(_10973_),
    .Y(_10984_));
 sky130_fd_sc_hd__nand2_2 _18948_ (.A(iX[1]),
    .B(iY[2]),
    .Y(_10995_));
 sky130_fd_sc_hd__xnor2_2 _18949_ (.A(_10984_),
    .B(_10995_),
    .Y(_11006_));
 sky130_fd_sc_hd__o21ba_2 _18950_ (.A1(_10875_),
    .A2(_10897_),
    .B1_N(_10864_),
    .X(_11016_));
 sky130_fd_sc_hd__xnor2_2 _18951_ (.A(_11006_),
    .B(_11016_),
    .Y(_11027_));
 sky130_fd_sc_hd__nand3_2 _18952_ (.A(iX[0]),
    .B(iY[3]),
    .C(_11027_),
    .Y(_11038_));
 sky130_fd_sc_hd__a21o_2 _18953_ (.A1(iX[0]),
    .A2(iY[3]),
    .B1(_11027_),
    .X(_11049_));
 sky130_fd_sc_hd__nand2_2 _18954_ (.A(_11038_),
    .B(_11049_),
    .Y(_11060_));
 sky130_fd_sc_hd__nor2_2 _18955_ (.A(_10919_),
    .B(_11060_),
    .Y(_11071_));
 sky130_fd_sc_hd__and2_2 _18956_ (.A(_10919_),
    .B(_11060_),
    .X(_11082_));
 sky130_fd_sc_hd__or2_2 _18957_ (.A(_11071_),
    .B(_11082_),
    .X(_11093_));
 sky130_fd_sc_hd__inv_2 _18958_ (.A(_11093_),
    .Y(oO[3]));
 sky130_fd_sc_hd__or2b_2 _18959_ (.A(_11016_),
    .B_N(_11006_),
    .X(_11114_));
 sky130_fd_sc_hd__and4_2 _18960_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[3]),
    .D(iX[4]),
    .X(_11125_));
 sky130_fd_sc_hd__a22o_2 _18961_ (.A1(iY[1]),
    .A2(iX[3]),
    .B1(iX[4]),
    .B2(iY[0]),
    .X(_11136_));
 sky130_fd_sc_hd__and2b_2 _18962_ (.A_N(_11125_),
    .B(_11136_),
    .X(_11147_));
 sky130_fd_sc_hd__nand2_2 _18963_ (.A(iX[2]),
    .B(iY[2]),
    .Y(_11158_));
 sky130_fd_sc_hd__xnor2_2 _18964_ (.A(_11147_),
    .B(_11158_),
    .Y(_11169_));
 sky130_fd_sc_hd__a31o_2 _18965_ (.A1(iX[1]),
    .A2(iY[2]),
    .A3(_10984_),
    .B1(_10962_),
    .X(_11180_));
 sky130_fd_sc_hd__xor2_2 _18966_ (.A(_11169_),
    .B(_11180_),
    .X(_11190_));
 sky130_fd_sc_hd__a22o_2 _18967_ (.A1(iX[1]),
    .A2(iY[3]),
    .B1(iY[4]),
    .B2(iX[0]),
    .X(_11201_));
 sky130_fd_sc_hd__nand4_2 _18968_ (.A(iX[0]),
    .B(iX[1]),
    .C(iY[3]),
    .D(iY[4]),
    .Y(_11212_));
 sky130_fd_sc_hd__and2_2 _18969_ (.A(_11201_),
    .B(_11212_),
    .X(_11223_));
 sky130_fd_sc_hd__xnor2_2 _18970_ (.A(_11190_),
    .B(_11223_),
    .Y(_11234_));
 sky130_fd_sc_hd__a21o_2 _18971_ (.A1(_11114_),
    .A2(_11038_),
    .B1(_11234_),
    .X(_11245_));
 sky130_fd_sc_hd__nand3_2 _18972_ (.A(_11114_),
    .B(_11038_),
    .C(_11234_),
    .Y(_11256_));
 sky130_fd_sc_hd__and2_2 _18973_ (.A(_11245_),
    .B(_11256_),
    .X(_11267_));
 sky130_fd_sc_hd__and2_2 _18974_ (.A(_11071_),
    .B(_11267_),
    .X(_11278_));
 sky130_fd_sc_hd__nor2_2 _18975_ (.A(_11071_),
    .B(_11267_),
    .Y(_11289_));
 sky130_fd_sc_hd__or2_2 _18976_ (.A(_11278_),
    .B(_11289_),
    .X(_11300_));
 sky130_fd_sc_hd__inv_2 _18977_ (.A(_11300_),
    .Y(oO[4]));
 sky130_fd_sc_hd__and4_2 _18978_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[4]),
    .D(iX[5]),
    .X(_11321_));
 sky130_fd_sc_hd__a22oi_2 _18979_ (.A1(iY[1]),
    .A2(iX[4]),
    .B1(iX[5]),
    .B2(iY[0]),
    .Y(_11332_));
 sky130_fd_sc_hd__nand2_2 _18980_ (.A(iY[2]),
    .B(iX[3]),
    .Y(_11343_));
 sky130_fd_sc_hd__or3_2 _18981_ (.A(_11321_),
    .B(_11332_),
    .C(_11343_),
    .X(_11354_));
 sky130_fd_sc_hd__o21ai_2 _18982_ (.A1(_11321_),
    .A2(_11332_),
    .B1(_11343_),
    .Y(_11365_));
 sky130_fd_sc_hd__a31o_2 _18983_ (.A1(iX[2]),
    .A2(iY[2]),
    .A3(_11136_),
    .B1(_11125_),
    .X(_11376_));
 sky130_fd_sc_hd__and3_2 _18984_ (.A(_11354_),
    .B(_11365_),
    .C(_11376_),
    .X(_11387_));
 sky130_fd_sc_hd__a21o_2 _18985_ (.A1(_11354_),
    .A2(_11365_),
    .B1(_11376_),
    .X(_11398_));
 sky130_fd_sc_hd__and2b_2 _18986_ (.A_N(_11387_),
    .B(_11398_),
    .X(_11409_));
 sky130_fd_sc_hd__and4_2 _18987_ (.A(iX[1]),
    .B(iX[2]),
    .C(iY[3]),
    .D(iY[4]),
    .X(_11420_));
 sky130_fd_sc_hd__a22oi_2 _18988_ (.A1(iX[2]),
    .A2(iY[3]),
    .B1(iY[4]),
    .B2(iX[1]),
    .Y(_11431_));
 sky130_fd_sc_hd__or2_2 _18989_ (.A(_11420_),
    .B(_11431_),
    .X(_11442_));
 sky130_fd_sc_hd__nand2_2 _18990_ (.A(iX[0]),
    .B(iY[5]),
    .Y(_11453_));
 sky130_fd_sc_hd__xor2_2 _18991_ (.A(_11442_),
    .B(_11453_),
    .X(_11464_));
 sky130_fd_sc_hd__xnor2_2 _18992_ (.A(_11409_),
    .B(_11464_),
    .Y(_11475_));
 sky130_fd_sc_hd__a22oi_2 _18993_ (.A1(_11169_),
    .A2(_11180_),
    .B1(_11190_),
    .B2(_11223_),
    .Y(_11486_));
 sky130_fd_sc_hd__xnor2_2 _18994_ (.A(_11475_),
    .B(_11486_),
    .Y(_11497_));
 sky130_fd_sc_hd__xnor2_2 _18995_ (.A(_11212_),
    .B(_11497_),
    .Y(_11508_));
 sky130_fd_sc_hd__xnor2_2 _18996_ (.A(_11245_),
    .B(_11508_),
    .Y(_11519_));
 sky130_fd_sc_hd__xnor2_2 _18997_ (.A(_11278_),
    .B(_11519_),
    .Y(oO[5]));
 sky130_fd_sc_hd__inv_2 _18998_ (.A(_11519_),
    .Y(_11540_));
 sky130_fd_sc_hd__nand2_2 _18999_ (.A(_11278_),
    .B(_11540_),
    .Y(_11551_));
 sky130_fd_sc_hd__and4_2 _19000_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[5]),
    .D(iX[6]),
    .X(_11562_));
 sky130_fd_sc_hd__a22oi_2 _19001_ (.A1(iY[1]),
    .A2(iX[5]),
    .B1(iX[6]),
    .B2(iY[0]),
    .Y(_11573_));
 sky130_fd_sc_hd__nand2_2 _19002_ (.A(iY[2]),
    .B(iX[4]),
    .Y(_11584_));
 sky130_fd_sc_hd__or3_2 _19003_ (.A(_11562_),
    .B(_11573_),
    .C(_11584_),
    .X(_11595_));
 sky130_fd_sc_hd__o21ai_2 _19004_ (.A1(_11562_),
    .A2(_11573_),
    .B1(_11584_),
    .Y(_11605_));
 sky130_fd_sc_hd__o21bai_2 _19005_ (.A1(_11332_),
    .A2(_11343_),
    .B1_N(_11321_),
    .Y(_11616_));
 sky130_fd_sc_hd__nand3_2 _19006_ (.A(_11595_),
    .B(_11605_),
    .C(_11616_),
    .Y(_11627_));
 sky130_fd_sc_hd__a21o_2 _19007_ (.A1(_11595_),
    .A2(_11605_),
    .B1(_11616_),
    .X(_11638_));
 sky130_fd_sc_hd__and4_2 _19008_ (.A(iX[2]),
    .B(iX[3]),
    .C(iY[3]),
    .D(iY[4]),
    .X(_11649_));
 sky130_fd_sc_hd__a22oi_2 _19009_ (.A1(iX[3]),
    .A2(iY[3]),
    .B1(iY[4]),
    .B2(iX[2]),
    .Y(_11660_));
 sky130_fd_sc_hd__nor2_2 _19010_ (.A(_11649_),
    .B(_11660_),
    .Y(_11671_));
 sky130_fd_sc_hd__nand2_2 _19011_ (.A(iX[1]),
    .B(iY[5]),
    .Y(_11682_));
 sky130_fd_sc_hd__xnor2_2 _19012_ (.A(_11671_),
    .B(_11682_),
    .Y(_11693_));
 sky130_fd_sc_hd__nand3_2 _19013_ (.A(_11627_),
    .B(_11638_),
    .C(_11693_),
    .Y(_11704_));
 sky130_fd_sc_hd__a21o_2 _19014_ (.A1(_11627_),
    .A2(_11638_),
    .B1(_11693_),
    .X(_11715_));
 sky130_fd_sc_hd__a21o_2 _19015_ (.A1(_11398_),
    .A2(_11464_),
    .B1(_11387_),
    .X(_11726_));
 sky130_fd_sc_hd__nand3_2 _19016_ (.A(_11704_),
    .B(_11715_),
    .C(_11726_),
    .Y(_11737_));
 sky130_fd_sc_hd__a21o_2 _19017_ (.A1(_11704_),
    .A2(_11715_),
    .B1(_11726_),
    .X(_11748_));
 sky130_fd_sc_hd__o21bai_2 _19018_ (.A1(_11431_),
    .A2(_11453_),
    .B1_N(_11420_),
    .Y(_11759_));
 sky130_fd_sc_hd__nand2_2 _19019_ (.A(iX[0]),
    .B(iY[6]),
    .Y(_11770_));
 sky130_fd_sc_hd__xnor2_2 _19020_ (.A(_11759_),
    .B(_11770_),
    .Y(_11781_));
 sky130_fd_sc_hd__and3_2 _19021_ (.A(_11737_),
    .B(_11748_),
    .C(_11781_),
    .X(_11792_));
 sky130_fd_sc_hd__a21oi_2 _19022_ (.A1(_11737_),
    .A2(_11748_),
    .B1(_11781_),
    .Y(_11803_));
 sky130_fd_sc_hd__nor2_2 _19023_ (.A(_11792_),
    .B(_11803_),
    .Y(_11814_));
 sky130_fd_sc_hd__or2_2 _19024_ (.A(_11475_),
    .B(_11486_),
    .X(_11824_));
 sky130_fd_sc_hd__o21a_2 _19025_ (.A1(_11212_),
    .A2(_11497_),
    .B1(_11824_),
    .X(_11835_));
 sky130_fd_sc_hd__xor2_2 _19026_ (.A(_11814_),
    .B(_11835_),
    .X(_11846_));
 sky130_fd_sc_hd__or2_2 _19027_ (.A(_11551_),
    .B(_11846_),
    .X(_11857_));
 sky130_fd_sc_hd__inv_2 _19028_ (.A(_11857_),
    .Y(_11868_));
 sky130_fd_sc_hd__or2_2 _19029_ (.A(_11245_),
    .B(_11508_),
    .X(_11879_));
 sky130_fd_sc_hd__nor2_2 _19030_ (.A(_11879_),
    .B(_11846_),
    .Y(_11890_));
 sky130_fd_sc_hd__or2_2 _19031_ (.A(_11868_),
    .B(_11890_),
    .X(_11901_));
 sky130_fd_sc_hd__and3_2 _19032_ (.A(_11879_),
    .B(_11551_),
    .C(_11846_),
    .X(_11912_));
 sky130_fd_sc_hd__or2_2 _19033_ (.A(_11901_),
    .B(_11912_),
    .X(_11923_));
 sky130_fd_sc_hd__inv_2 _19034_ (.A(_11923_),
    .Y(oO[6]));
 sky130_fd_sc_hd__and2b_2 _19035_ (.A_N(_11835_),
    .B(_11814_),
    .X(_11944_));
 sky130_fd_sc_hd__and3_2 _19036_ (.A(iX[0]),
    .B(iY[6]),
    .C(_11759_),
    .X(_11955_));
 sky130_fd_sc_hd__and3_2 _19037_ (.A(_11704_),
    .B(_11715_),
    .C(_11726_),
    .X(_11966_));
 sky130_fd_sc_hd__and4_2 _19038_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[6]),
    .D(iX[7]),
    .X(_11977_));
 sky130_fd_sc_hd__a22oi_2 _19039_ (.A1(iY[1]),
    .A2(iX[6]),
    .B1(iX[7]),
    .B2(iY[0]),
    .Y(_11988_));
 sky130_fd_sc_hd__nand2_2 _19040_ (.A(iY[2]),
    .B(iX[5]),
    .Y(_11999_));
 sky130_fd_sc_hd__or3_2 _19041_ (.A(_11977_),
    .B(_11988_),
    .C(_11999_),
    .X(_12010_));
 sky130_fd_sc_hd__o21ai_2 _19042_ (.A1(_11977_),
    .A2(_11988_),
    .B1(_11999_),
    .Y(_12021_));
 sky130_fd_sc_hd__o21bai_2 _19043_ (.A1(_11573_),
    .A2(_11584_),
    .B1_N(_11562_),
    .Y(_12032_));
 sky130_fd_sc_hd__nand3_2 _19044_ (.A(_12010_),
    .B(_12021_),
    .C(_12032_),
    .Y(_12043_));
 sky130_fd_sc_hd__a21o_2 _19045_ (.A1(_12010_),
    .A2(_12021_),
    .B1(_12032_),
    .X(_12053_));
 sky130_fd_sc_hd__and4_2 _19046_ (.A(iX[3]),
    .B(iY[3]),
    .C(iX[4]),
    .D(iY[4]),
    .X(_12064_));
 sky130_fd_sc_hd__a22o_2 _19047_ (.A1(iY[3]),
    .A2(iX[4]),
    .B1(iY[4]),
    .B2(iX[3]),
    .X(_12075_));
 sky130_fd_sc_hd__and2b_2 _19048_ (.A_N(_12064_),
    .B(_12075_),
    .X(_12086_));
 sky130_fd_sc_hd__nand2_2 _19049_ (.A(iX[2]),
    .B(iY[5]),
    .Y(_12097_));
 sky130_fd_sc_hd__xnor2_2 _19050_ (.A(_12086_),
    .B(_12097_),
    .Y(_12108_));
 sky130_fd_sc_hd__nand3_2 _19051_ (.A(_12043_),
    .B(_12053_),
    .C(_12108_),
    .Y(_12119_));
 sky130_fd_sc_hd__a21o_2 _19052_ (.A1(_12043_),
    .A2(_12053_),
    .B1(_12108_),
    .X(_12130_));
 sky130_fd_sc_hd__a21bo_2 _19053_ (.A1(_11638_),
    .A2(_11693_),
    .B1_N(_11627_),
    .X(_12141_));
 sky130_fd_sc_hd__nand3_2 _19054_ (.A(_12119_),
    .B(_12130_),
    .C(_12141_),
    .Y(_12152_));
 sky130_fd_sc_hd__a21o_2 _19055_ (.A1(_12119_),
    .A2(_12130_),
    .B1(_12141_),
    .X(_12163_));
 sky130_fd_sc_hd__a31o_2 _19056_ (.A1(iX[1]),
    .A2(iY[5]),
    .A3(_11671_),
    .B1(_11649_),
    .X(_12174_));
 sky130_fd_sc_hd__and4_2 _19057_ (.A(iX[0]),
    .B(iX[1]),
    .C(iY[6]),
    .D(iY[7]),
    .X(_12185_));
 sky130_fd_sc_hd__a22oi_2 _19058_ (.A1(iX[1]),
    .A2(iY[6]),
    .B1(iY[7]),
    .B2(iX[0]),
    .Y(_12196_));
 sky130_fd_sc_hd__or2_2 _19059_ (.A(_12185_),
    .B(_12196_),
    .X(_12207_));
 sky130_fd_sc_hd__xnor2_2 _19060_ (.A(_12174_),
    .B(_12207_),
    .Y(_12218_));
 sky130_fd_sc_hd__nand3_2 _19061_ (.A(_12152_),
    .B(_12163_),
    .C(_12218_),
    .Y(_12229_));
 sky130_fd_sc_hd__a21o_2 _19062_ (.A1(_12152_),
    .A2(_12163_),
    .B1(_12218_),
    .X(_12240_));
 sky130_fd_sc_hd__o211ai_2 _19063_ (.A1(_11966_),
    .A2(_11792_),
    .B1(_12229_),
    .C1(_12240_),
    .Y(_12251_));
 sky130_fd_sc_hd__a211o_2 _19064_ (.A1(_12229_),
    .A2(_12240_),
    .B1(_11966_),
    .C1(_11792_),
    .X(_12262_));
 sky130_fd_sc_hd__nand3_2 _19065_ (.A(_11955_),
    .B(_12251_),
    .C(_12262_),
    .Y(_12273_));
 sky130_fd_sc_hd__a21o_2 _19066_ (.A1(_12251_),
    .A2(_12262_),
    .B1(_11955_),
    .X(_12284_));
 sky130_fd_sc_hd__and3_2 _19067_ (.A(_11944_),
    .B(_12273_),
    .C(_12284_),
    .X(_12294_));
 sky130_fd_sc_hd__a21o_2 _19068_ (.A1(_12273_),
    .A2(_12284_),
    .B1(_11944_),
    .X(_12305_));
 sky130_fd_sc_hd__and2b_2 _19069_ (.A_N(_12294_),
    .B(_12305_),
    .X(_12316_));
 sky130_fd_sc_hd__xnor2_2 _19070_ (.A(_11901_),
    .B(_12316_),
    .Y(_12327_));
 sky130_fd_sc_hd__inv_2 _19071_ (.A(_12327_),
    .Y(oO[7]));
 sky130_fd_sc_hd__and2_2 _19072_ (.A(_11868_),
    .B(_12316_),
    .X(_12348_));
 sky130_fd_sc_hd__and2b_2 _19073_ (.A_N(_12207_),
    .B(_12174_),
    .X(_12359_));
 sky130_fd_sc_hd__and4_2 _19074_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[7]),
    .D(iX[8]),
    .X(_12370_));
 sky130_fd_sc_hd__a22oi_2 _19075_ (.A1(iY[1]),
    .A2(iX[7]),
    .B1(iX[8]),
    .B2(iY[0]),
    .Y(_12381_));
 sky130_fd_sc_hd__nand2_2 _19076_ (.A(iY[2]),
    .B(iX[6]),
    .Y(_12392_));
 sky130_fd_sc_hd__or3_2 _19077_ (.A(_12370_),
    .B(_12381_),
    .C(_12392_),
    .X(_12403_));
 sky130_fd_sc_hd__o21ai_2 _19078_ (.A1(_12370_),
    .A2(_12381_),
    .B1(_12392_),
    .Y(_12414_));
 sky130_fd_sc_hd__o21bai_2 _19079_ (.A1(_11988_),
    .A2(_11999_),
    .B1_N(_11977_),
    .Y(_12425_));
 sky130_fd_sc_hd__nand3_2 _19080_ (.A(_12403_),
    .B(_12414_),
    .C(_12425_),
    .Y(_12436_));
 sky130_fd_sc_hd__a21o_2 _19081_ (.A1(_12403_),
    .A2(_12414_),
    .B1(_12425_),
    .X(_12447_));
 sky130_fd_sc_hd__and4_2 _19082_ (.A(iY[3]),
    .B(iX[4]),
    .C(iY[4]),
    .D(iX[5]),
    .X(_12458_));
 sky130_fd_sc_hd__a22oi_2 _19083_ (.A1(iX[4]),
    .A2(iY[4]),
    .B1(iX[5]),
    .B2(iY[3]),
    .Y(_12469_));
 sky130_fd_sc_hd__nor2_2 _19084_ (.A(_12458_),
    .B(_12469_),
    .Y(_12480_));
 sky130_fd_sc_hd__nand2_2 _19085_ (.A(iX[3]),
    .B(iY[5]),
    .Y(_12491_));
 sky130_fd_sc_hd__xnor2_2 _19086_ (.A(_12480_),
    .B(_12491_),
    .Y(_12502_));
 sky130_fd_sc_hd__nand3_2 _19087_ (.A(_12436_),
    .B(_12447_),
    .C(_12502_),
    .Y(_12513_));
 sky130_fd_sc_hd__a21o_2 _19088_ (.A1(_12436_),
    .A2(_12447_),
    .B1(_12502_),
    .X(_12524_));
 sky130_fd_sc_hd__a21bo_2 _19089_ (.A1(_12053_),
    .A2(_12108_),
    .B1_N(_12043_),
    .X(_12535_));
 sky130_fd_sc_hd__and3_2 _19090_ (.A(_12513_),
    .B(_12524_),
    .C(_12535_),
    .X(_12545_));
 sky130_fd_sc_hd__a21oi_2 _19091_ (.A1(_12513_),
    .A2(_12524_),
    .B1(_12535_),
    .Y(_12556_));
 sky130_fd_sc_hd__a31o_2 _19092_ (.A1(iX[2]),
    .A2(iY[5]),
    .A3(_12075_),
    .B1(_12064_),
    .X(_12567_));
 sky130_fd_sc_hd__and4_2 _19093_ (.A(iX[1]),
    .B(iX[2]),
    .C(iY[6]),
    .D(iY[7]),
    .X(_12578_));
 sky130_fd_sc_hd__a22oi_2 _19094_ (.A1(iX[2]),
    .A2(iY[6]),
    .B1(iY[7]),
    .B2(iX[1]),
    .Y(_12589_));
 sky130_fd_sc_hd__nor2_2 _19095_ (.A(_12578_),
    .B(_12589_),
    .Y(_12600_));
 sky130_fd_sc_hd__nand2_2 _19096_ (.A(iX[0]),
    .B(iY[8]),
    .Y(_12611_));
 sky130_fd_sc_hd__xnor2_2 _19097_ (.A(_12600_),
    .B(_12611_),
    .Y(_12622_));
 sky130_fd_sc_hd__xor2_2 _19098_ (.A(_12567_),
    .B(_12622_),
    .X(_12633_));
 sky130_fd_sc_hd__xnor2_2 _19099_ (.A(_12185_),
    .B(_12633_),
    .Y(_12644_));
 sky130_fd_sc_hd__nor3_2 _19100_ (.A(_12545_),
    .B(_12556_),
    .C(_12644_),
    .Y(_12655_));
 sky130_fd_sc_hd__o21a_2 _19101_ (.A1(_12545_),
    .A2(_12556_),
    .B1(_12644_),
    .X(_12666_));
 sky130_fd_sc_hd__a211o_2 _19102_ (.A1(_12152_),
    .A2(_12229_),
    .B1(_12655_),
    .C1(_12666_),
    .X(_12677_));
 sky130_fd_sc_hd__o211ai_2 _19103_ (.A1(_12655_),
    .A2(_12666_),
    .B1(_12152_),
    .C1(_12229_),
    .Y(_12688_));
 sky130_fd_sc_hd__and3_2 _19104_ (.A(_12359_),
    .B(_12677_),
    .C(_12688_),
    .X(_12699_));
 sky130_fd_sc_hd__a21oi_2 _19105_ (.A1(_12677_),
    .A2(_12688_),
    .B1(_12359_),
    .Y(_12710_));
 sky130_fd_sc_hd__a211o_2 _19106_ (.A1(_12251_),
    .A2(_12273_),
    .B1(_12699_),
    .C1(_12710_),
    .X(_12721_));
 sky130_fd_sc_hd__o211ai_2 _19107_ (.A1(_12699_),
    .A2(_12710_),
    .B1(_12251_),
    .C1(_12273_),
    .Y(_12732_));
 sky130_fd_sc_hd__nand2_2 _19108_ (.A(_12721_),
    .B(_12732_),
    .Y(_12743_));
 sky130_fd_sc_hd__a21oi_2 _19109_ (.A1(_11890_),
    .A2(_12305_),
    .B1(_12294_),
    .Y(_12754_));
 sky130_fd_sc_hd__xnor2_2 _19110_ (.A(_12743_),
    .B(_12754_),
    .Y(_12765_));
 sky130_fd_sc_hd__xor2_2 _19111_ (.A(_12348_),
    .B(_12765_),
    .X(_12776_));
 sky130_fd_sc_hd__inv_2 _19112_ (.A(_12776_),
    .Y(oO[8]));
 sky130_fd_sc_hd__a211oi_2 _19113_ (.A1(_12251_),
    .A2(_12273_),
    .B1(_12699_),
    .C1(_12710_),
    .Y(_12797_));
 sky130_fd_sc_hd__a211oi_2 _19114_ (.A1(_12152_),
    .A2(_12229_),
    .B1(_12655_),
    .C1(_12666_),
    .Y(_12807_));
 sky130_fd_sc_hd__and4_2 _19115_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[8]),
    .D(iX[9]),
    .X(_12818_));
 sky130_fd_sc_hd__a22oi_2 _19116_ (.A1(iY[1]),
    .A2(iX[8]),
    .B1(iX[9]),
    .B2(iY[0]),
    .Y(_12829_));
 sky130_fd_sc_hd__nand2_2 _19117_ (.A(iY[2]),
    .B(iX[7]),
    .Y(_12840_));
 sky130_fd_sc_hd__or3_2 _19118_ (.A(_12818_),
    .B(_12829_),
    .C(_12840_),
    .X(_12851_));
 sky130_fd_sc_hd__o21ai_2 _19119_ (.A1(_12818_),
    .A2(_12829_),
    .B1(_12840_),
    .Y(_12862_));
 sky130_fd_sc_hd__o21bai_2 _19120_ (.A1(_12381_),
    .A2(_12392_),
    .B1_N(_12370_),
    .Y(_12873_));
 sky130_fd_sc_hd__nand3_2 _19121_ (.A(_12851_),
    .B(_12862_),
    .C(_12873_),
    .Y(_12884_));
 sky130_fd_sc_hd__a21o_2 _19122_ (.A1(_12851_),
    .A2(_12862_),
    .B1(_12873_),
    .X(_12895_));
 sky130_fd_sc_hd__and4_2 _19123_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[5]),
    .D(iX[6]),
    .X(_12906_));
 sky130_fd_sc_hd__a22oi_2 _19124_ (.A1(iY[4]),
    .A2(iX[5]),
    .B1(iX[6]),
    .B2(iY[3]),
    .Y(_12917_));
 sky130_fd_sc_hd__nor2_2 _19125_ (.A(_12906_),
    .B(_12917_),
    .Y(_12928_));
 sky130_fd_sc_hd__nand2_2 _19126_ (.A(iX[4]),
    .B(iY[5]),
    .Y(_12939_));
 sky130_fd_sc_hd__xnor2_2 _19127_ (.A(_12928_),
    .B(_12939_),
    .Y(_12950_));
 sky130_fd_sc_hd__nand3_2 _19128_ (.A(_12884_),
    .B(_12895_),
    .C(_12950_),
    .Y(_12961_));
 sky130_fd_sc_hd__a21o_2 _19129_ (.A1(_12884_),
    .A2(_12895_),
    .B1(_12950_),
    .X(_12972_));
 sky130_fd_sc_hd__a21bo_2 _19130_ (.A1(_12447_),
    .A2(_12502_),
    .B1_N(_12436_),
    .X(_12983_));
 sky130_fd_sc_hd__nand3_2 _19131_ (.A(_12961_),
    .B(_12972_),
    .C(_12983_),
    .Y(_12994_));
 sky130_fd_sc_hd__a21o_2 _19132_ (.A1(_12961_),
    .A2(_12972_),
    .B1(_12983_),
    .X(_13005_));
 sky130_fd_sc_hd__o21ba_2 _19133_ (.A1(_12589_),
    .A2(_12611_),
    .B1_N(_12578_),
    .X(_13016_));
 sky130_fd_sc_hd__o21ba_2 _19134_ (.A1(_12469_),
    .A2(_12491_),
    .B1_N(_12458_),
    .X(_13027_));
 sky130_fd_sc_hd__and4_2 _19135_ (.A(iX[2]),
    .B(iX[3]),
    .C(iY[6]),
    .D(iY[7]),
    .X(_13038_));
 sky130_fd_sc_hd__a22oi_2 _19136_ (.A1(iX[3]),
    .A2(iY[6]),
    .B1(iY[7]),
    .B2(iX[2]),
    .Y(_13049_));
 sky130_fd_sc_hd__nor2_2 _19137_ (.A(_13038_),
    .B(_13049_),
    .Y(_13060_));
 sky130_fd_sc_hd__nand2_2 _19138_ (.A(iX[1]),
    .B(iY[8]),
    .Y(_13070_));
 sky130_fd_sc_hd__xnor2_2 _19139_ (.A(_13060_),
    .B(_13070_),
    .Y(_13081_));
 sky130_fd_sc_hd__xnor2_2 _19140_ (.A(_13027_),
    .B(_13081_),
    .Y(_13092_));
 sky130_fd_sc_hd__xnor2_2 _19141_ (.A(_13016_),
    .B(_13092_),
    .Y(_13103_));
 sky130_fd_sc_hd__nand3_2 _19142_ (.A(_12994_),
    .B(_13005_),
    .C(_13103_),
    .Y(_13114_));
 sky130_fd_sc_hd__a21o_2 _19143_ (.A1(_12994_),
    .A2(_13005_),
    .B1(_13103_),
    .X(_13125_));
 sky130_fd_sc_hd__o211ai_2 _19144_ (.A1(_12545_),
    .A2(_12655_),
    .B1(_13114_),
    .C1(_13125_),
    .Y(_13136_));
 sky130_fd_sc_hd__a211o_2 _19145_ (.A1(_13114_),
    .A2(_13125_),
    .B1(_12545_),
    .C1(_12655_),
    .X(_13147_));
 sky130_fd_sc_hd__and2_2 _19146_ (.A(_12567_),
    .B(_12622_),
    .X(_13158_));
 sky130_fd_sc_hd__and2_2 _19147_ (.A(_12185_),
    .B(_12633_),
    .X(_13169_));
 sky130_fd_sc_hd__o211a_2 _19148_ (.A1(_13158_),
    .A2(_13169_),
    .B1(iX[0]),
    .C1(iY[9]),
    .X(_13180_));
 sky130_fd_sc_hd__a211oi_2 _19149_ (.A1(iX[0]),
    .A2(iY[9]),
    .B1(_13158_),
    .C1(_13169_),
    .Y(_13191_));
 sky130_fd_sc_hd__nor2_2 _19150_ (.A(_13180_),
    .B(_13191_),
    .Y(_13202_));
 sky130_fd_sc_hd__nand3_2 _19151_ (.A(_13136_),
    .B(_13147_),
    .C(_13202_),
    .Y(_13213_));
 sky130_fd_sc_hd__a21o_2 _19152_ (.A1(_13136_),
    .A2(_13147_),
    .B1(_13202_),
    .X(_13224_));
 sky130_fd_sc_hd__o211ai_2 _19153_ (.A1(_12807_),
    .A2(_12699_),
    .B1(_13213_),
    .C1(_13224_),
    .Y(_13235_));
 sky130_fd_sc_hd__a211o_2 _19154_ (.A1(_13213_),
    .A2(_13224_),
    .B1(_12807_),
    .C1(_12699_),
    .X(_13246_));
 sky130_fd_sc_hd__and3_2 _19155_ (.A(_12797_),
    .B(_13235_),
    .C(_13246_),
    .X(_13257_));
 sky130_fd_sc_hd__a21o_2 _19156_ (.A1(_13235_),
    .A2(_13246_),
    .B1(_12797_),
    .X(_13268_));
 sky130_fd_sc_hd__and2b_2 _19157_ (.A_N(_13257_),
    .B(_13268_),
    .X(_13279_));
 sky130_fd_sc_hd__and3_2 _19158_ (.A(_12294_),
    .B(_12721_),
    .C(_12732_),
    .X(_13290_));
 sky130_fd_sc_hd__and4bb_2 _19159_ (.A_N(_12294_),
    .B_N(_12743_),
    .C(_12305_),
    .D(_11890_),
    .X(_13301_));
 sky130_fd_sc_hd__or4b_2 _19160_ (.A(_11857_),
    .B(_12294_),
    .C(_12765_),
    .D_N(_12305_),
    .X(_13312_));
 sky130_fd_sc_hd__or3b_2 _19161_ (.A(_13290_),
    .B(_13301_),
    .C_N(_13312_),
    .X(_13323_));
 sky130_fd_sc_hd__xor2_2 _19162_ (.A(_13279_),
    .B(_13323_),
    .X(oO[9]));
 sky130_fd_sc_hd__o211a_2 _19163_ (.A1(_12545_),
    .A2(_12655_),
    .B1(_13114_),
    .C1(_13125_),
    .X(_13344_));
 sky130_fd_sc_hd__and3_2 _19164_ (.A(_13136_),
    .B(_13147_),
    .C(_13202_),
    .X(_13354_));
 sky130_fd_sc_hd__nand2_2 _19165_ (.A(iY[2]),
    .B(iX[8]),
    .Y(_13365_));
 sky130_fd_sc_hd__a22o_2 _19166_ (.A1(iY[1]),
    .A2(iX[9]),
    .B1(iX[10]),
    .B2(iY[0]),
    .X(_13376_));
 sky130_fd_sc_hd__nand4_2 _19167_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[9]),
    .D(iX[10]),
    .Y(_13387_));
 sky130_fd_sc_hd__nand3b_2 _19168_ (.A_N(_13365_),
    .B(_13376_),
    .C(_13387_),
    .Y(_13398_));
 sky130_fd_sc_hd__a21bo_2 _19169_ (.A1(_13387_),
    .A2(_13376_),
    .B1_N(_13365_),
    .X(_13409_));
 sky130_fd_sc_hd__o21bai_2 _19170_ (.A1(_12829_),
    .A2(_12840_),
    .B1_N(_12818_),
    .Y(_13420_));
 sky130_fd_sc_hd__nand3_2 _19171_ (.A(_13398_),
    .B(_13409_),
    .C(_13420_),
    .Y(_13431_));
 sky130_fd_sc_hd__a21o_2 _19172_ (.A1(_13398_),
    .A2(_13409_),
    .B1(_13420_),
    .X(_13442_));
 sky130_fd_sc_hd__and4_2 _19173_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[6]),
    .D(iX[7]),
    .X(_13453_));
 sky130_fd_sc_hd__a22oi_2 _19174_ (.A1(iY[4]),
    .A2(iX[6]),
    .B1(iX[7]),
    .B2(iY[3]),
    .Y(_13464_));
 sky130_fd_sc_hd__nor2_2 _19175_ (.A(_13453_),
    .B(_13464_),
    .Y(_13475_));
 sky130_fd_sc_hd__nand2_2 _19176_ (.A(iX[5]),
    .B(iY[5]),
    .Y(_13486_));
 sky130_fd_sc_hd__xnor2_2 _19177_ (.A(_13475_),
    .B(_13486_),
    .Y(_13497_));
 sky130_fd_sc_hd__nand3_2 _19178_ (.A(_13431_),
    .B(_13442_),
    .C(_13497_),
    .Y(_13508_));
 sky130_fd_sc_hd__a21o_2 _19179_ (.A1(_13431_),
    .A2(_13442_),
    .B1(_13497_),
    .X(_13519_));
 sky130_fd_sc_hd__a21bo_2 _19180_ (.A1(_12895_),
    .A2(_12950_),
    .B1_N(_12884_),
    .X(_13530_));
 sky130_fd_sc_hd__nand3_2 _19181_ (.A(_13508_),
    .B(_13519_),
    .C(_13530_),
    .Y(_13541_));
 sky130_fd_sc_hd__a21o_2 _19182_ (.A1(_13508_),
    .A2(_13519_),
    .B1(_13530_),
    .X(_13552_));
 sky130_fd_sc_hd__o21ba_2 _19183_ (.A1(_13049_),
    .A2(_13070_),
    .B1_N(_13038_),
    .X(_13563_));
 sky130_fd_sc_hd__o21ba_2 _19184_ (.A1(_12917_),
    .A2(_12939_),
    .B1_N(_12906_),
    .X(_13574_));
 sky130_fd_sc_hd__and4_2 _19185_ (.A(iX[3]),
    .B(iX[4]),
    .C(iY[6]),
    .D(iY[7]),
    .X(_13585_));
 sky130_fd_sc_hd__a22oi_2 _19186_ (.A1(iX[4]),
    .A2(iY[6]),
    .B1(iY[7]),
    .B2(iX[3]),
    .Y(_13596_));
 sky130_fd_sc_hd__nor2_2 _19187_ (.A(_13585_),
    .B(_13596_),
    .Y(_13607_));
 sky130_fd_sc_hd__nand2_2 _19188_ (.A(iX[2]),
    .B(iY[8]),
    .Y(_13618_));
 sky130_fd_sc_hd__xnor2_2 _19189_ (.A(_13607_),
    .B(_13618_),
    .Y(_13629_));
 sky130_fd_sc_hd__xnor2_2 _19190_ (.A(_13574_),
    .B(_13629_),
    .Y(_13639_));
 sky130_fd_sc_hd__xnor2_2 _19191_ (.A(_13563_),
    .B(_13639_),
    .Y(_13650_));
 sky130_fd_sc_hd__and3_2 _19192_ (.A(_13541_),
    .B(_13552_),
    .C(_13650_),
    .X(_13661_));
 sky130_fd_sc_hd__a21oi_2 _19193_ (.A1(_13541_),
    .A2(_13552_),
    .B1(_13650_),
    .Y(_13672_));
 sky130_fd_sc_hd__a211o_2 _19194_ (.A1(_12994_),
    .A2(_13114_),
    .B1(_13661_),
    .C1(_13672_),
    .X(_13683_));
 sky130_fd_sc_hd__o211ai_2 _19195_ (.A1(_13661_),
    .A2(_13672_),
    .B1(_12994_),
    .C1(_13114_),
    .Y(_13694_));
 sky130_fd_sc_hd__or2b_2 _19196_ (.A(_13027_),
    .B_N(_13081_),
    .X(_13705_));
 sky130_fd_sc_hd__or2b_2 _19197_ (.A(_13016_),
    .B_N(_13092_),
    .X(_13716_));
 sky130_fd_sc_hd__a22oi_2 _19198_ (.A1(iX[1]),
    .A2(iY[9]),
    .B1(iY[10]),
    .B2(iX[0]),
    .Y(_13727_));
 sky130_fd_sc_hd__and4_2 _19199_ (.A(iX[0]),
    .B(iX[1]),
    .C(iY[9]),
    .D(iY[10]),
    .X(_13738_));
 sky130_fd_sc_hd__or2_2 _19200_ (.A(_13727_),
    .B(_13738_),
    .X(_13749_));
 sky130_fd_sc_hd__a21oi_2 _19201_ (.A1(_13705_),
    .A2(_13716_),
    .B1(_13749_),
    .Y(_13760_));
 sky130_fd_sc_hd__and3_2 _19202_ (.A(_13705_),
    .B(_13716_),
    .C(_13749_),
    .X(_13771_));
 sky130_fd_sc_hd__nor2_2 _19203_ (.A(_13760_),
    .B(_13771_),
    .Y(_13782_));
 sky130_fd_sc_hd__nand3_2 _19204_ (.A(_13683_),
    .B(_13694_),
    .C(_13782_),
    .Y(_13793_));
 sky130_fd_sc_hd__a21o_2 _19205_ (.A1(_13683_),
    .A2(_13694_),
    .B1(_13782_),
    .X(_13804_));
 sky130_fd_sc_hd__o211ai_2 _19206_ (.A1(_13344_),
    .A2(_13354_),
    .B1(_13793_),
    .C1(_13804_),
    .Y(_13815_));
 sky130_fd_sc_hd__a211o_2 _19207_ (.A1(_13793_),
    .A2(_13804_),
    .B1(_13344_),
    .C1(_13354_),
    .X(_13826_));
 sky130_fd_sc_hd__and3_2 _19208_ (.A(_13180_),
    .B(_13815_),
    .C(_13826_),
    .X(_13837_));
 sky130_fd_sc_hd__a21oi_2 _19209_ (.A1(_13815_),
    .A2(_13826_),
    .B1(_13180_),
    .Y(_13848_));
 sky130_fd_sc_hd__or3_2 _19210_ (.A(_13235_),
    .B(_13837_),
    .C(_13848_),
    .X(_13859_));
 sky130_fd_sc_hd__o21ai_2 _19211_ (.A1(_13837_),
    .A2(_13848_),
    .B1(_13235_),
    .Y(_13870_));
 sky130_fd_sc_hd__a21oi_2 _19212_ (.A1(_13290_),
    .A2(_13268_),
    .B1(_13257_),
    .Y(_13881_));
 sky130_fd_sc_hd__and3_2 _19213_ (.A(_13859_),
    .B(_13870_),
    .C(_13881_),
    .X(_13892_));
 sky130_fd_sc_hd__a21oi_2 _19214_ (.A1(_13859_),
    .A2(_13870_),
    .B1(_13881_),
    .Y(_13903_));
 sky130_fd_sc_hd__and2_2 _19215_ (.A(_13301_),
    .B(_13279_),
    .X(_13914_));
 sky130_fd_sc_hd__o21a_2 _19216_ (.A1(_13892_),
    .A2(_13903_),
    .B1(_13914_),
    .X(_13924_));
 sky130_fd_sc_hd__nor3_2 _19217_ (.A(_13914_),
    .B(_13892_),
    .C(_13903_),
    .Y(_13935_));
 sky130_fd_sc_hd__nor2_2 _19218_ (.A(_13924_),
    .B(_13935_),
    .Y(_13946_));
 sky130_fd_sc_hd__or2b_2 _19219_ (.A(_13312_),
    .B_N(_13279_),
    .X(_13957_));
 sky130_fd_sc_hd__xnor2_2 _19220_ (.A(_13946_),
    .B(_13957_),
    .Y(oO[10]));
 sky130_fd_sc_hd__nand2_2 _19221_ (.A(_13290_),
    .B(_13279_),
    .Y(_13978_));
 sky130_fd_sc_hd__nand2_2 _19222_ (.A(_13859_),
    .B(_13870_),
    .Y(_13989_));
 sky130_fd_sc_hd__and4_2 _19223_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[10]),
    .D(iX[11]),
    .X(_14000_));
 sky130_fd_sc_hd__a22oi_2 _19224_ (.A1(iY[1]),
    .A2(iX[10]),
    .B1(iX[11]),
    .B2(iY[0]),
    .Y(_14011_));
 sky130_fd_sc_hd__nor2_2 _19225_ (.A(_14000_),
    .B(_14011_),
    .Y(_14022_));
 sky130_fd_sc_hd__nand2_2 _19226_ (.A(iY[2]),
    .B(iX[9]),
    .Y(_14033_));
 sky130_fd_sc_hd__xnor2_2 _19227_ (.A(_14022_),
    .B(_14033_),
    .Y(_14044_));
 sky130_fd_sc_hd__nand2_2 _19228_ (.A(_13387_),
    .B(_13398_),
    .Y(_14055_));
 sky130_fd_sc_hd__xor2_2 _19229_ (.A(_14044_),
    .B(_14055_),
    .X(_14066_));
 sky130_fd_sc_hd__and4_2 _19230_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[7]),
    .D(iX[8]),
    .X(_14077_));
 sky130_fd_sc_hd__a22oi_2 _19231_ (.A1(iY[4]),
    .A2(iX[7]),
    .B1(iX[8]),
    .B2(iY[3]),
    .Y(_14088_));
 sky130_fd_sc_hd__nor2_2 _19232_ (.A(_14077_),
    .B(_14088_),
    .Y(_14099_));
 sky130_fd_sc_hd__nand2_2 _19233_ (.A(iY[5]),
    .B(iX[6]),
    .Y(_14110_));
 sky130_fd_sc_hd__xnor2_2 _19234_ (.A(_14099_),
    .B(_14110_),
    .Y(_14121_));
 sky130_fd_sc_hd__xnor2_2 _19235_ (.A(_14066_),
    .B(_14121_),
    .Y(_14132_));
 sky130_fd_sc_hd__and2_2 _19236_ (.A(_13431_),
    .B(_13508_),
    .X(_14143_));
 sky130_fd_sc_hd__xor2_2 _19237_ (.A(_14132_),
    .B(_14143_),
    .X(_14154_));
 sky130_fd_sc_hd__o21ba_2 _19238_ (.A1(_13596_),
    .A2(_13618_),
    .B1_N(_13585_),
    .X(_14165_));
 sky130_fd_sc_hd__o21ba_2 _19239_ (.A1(_13464_),
    .A2(_13486_),
    .B1_N(_13453_),
    .X(_14176_));
 sky130_fd_sc_hd__and4_2 _19240_ (.A(iX[4]),
    .B(iX[5]),
    .C(iY[6]),
    .D(iY[7]),
    .X(_14187_));
 sky130_fd_sc_hd__a22oi_2 _19241_ (.A1(iX[5]),
    .A2(iY[6]),
    .B1(iY[7]),
    .B2(iX[4]),
    .Y(_14198_));
 sky130_fd_sc_hd__nor2_2 _19242_ (.A(_14187_),
    .B(_14198_),
    .Y(_14209_));
 sky130_fd_sc_hd__nand2_2 _19243_ (.A(iX[3]),
    .B(iY[8]),
    .Y(_14219_));
 sky130_fd_sc_hd__xnor2_2 _19244_ (.A(_14209_),
    .B(_14219_),
    .Y(_14230_));
 sky130_fd_sc_hd__xnor2_2 _19245_ (.A(_14176_),
    .B(_14230_),
    .Y(_14241_));
 sky130_fd_sc_hd__xnor2_2 _19246_ (.A(_14165_),
    .B(_14241_),
    .Y(_14252_));
 sky130_fd_sc_hd__xnor2_2 _19247_ (.A(_14154_),
    .B(_14252_),
    .Y(_14263_));
 sky130_fd_sc_hd__a31o_2 _19248_ (.A1(_13508_),
    .A2(_13519_),
    .A3(_13530_),
    .B1(_13661_),
    .X(_14274_));
 sky130_fd_sc_hd__xnor2_2 _19249_ (.A(_14263_),
    .B(_14274_),
    .Y(_14285_));
 sky130_fd_sc_hd__or2b_2 _19250_ (.A(_13574_),
    .B_N(_13629_),
    .X(_14296_));
 sky130_fd_sc_hd__or2b_2 _19251_ (.A(_13563_),
    .B_N(_13639_),
    .X(_14307_));
 sky130_fd_sc_hd__and4_2 _19252_ (.A(iX[1]),
    .B(iX[2]),
    .C(iY[9]),
    .D(iY[10]),
    .X(_14318_));
 sky130_fd_sc_hd__a22oi_2 _19253_ (.A1(iX[2]),
    .A2(iY[9]),
    .B1(iY[10]),
    .B2(iX[1]),
    .Y(_14329_));
 sky130_fd_sc_hd__nor2_2 _19254_ (.A(_14318_),
    .B(_14329_),
    .Y(_14340_));
 sky130_fd_sc_hd__nand2_2 _19255_ (.A(iX[0]),
    .B(iY[11]),
    .Y(_14351_));
 sky130_fd_sc_hd__xnor2_2 _19256_ (.A(_14340_),
    .B(_14351_),
    .Y(_14362_));
 sky130_fd_sc_hd__and2_2 _19257_ (.A(_13738_),
    .B(_14362_),
    .X(_14373_));
 sky130_fd_sc_hd__nor2_2 _19258_ (.A(_13738_),
    .B(_14362_),
    .Y(_14384_));
 sky130_fd_sc_hd__or2_2 _19259_ (.A(_14373_),
    .B(_14384_),
    .X(_14395_));
 sky130_fd_sc_hd__a21oi_2 _19260_ (.A1(_14296_),
    .A2(_14307_),
    .B1(_14395_),
    .Y(_14406_));
 sky130_fd_sc_hd__and3_2 _19261_ (.A(_14296_),
    .B(_14307_),
    .C(_14395_),
    .X(_14417_));
 sky130_fd_sc_hd__nor2_2 _19262_ (.A(_14406_),
    .B(_14417_),
    .Y(_14428_));
 sky130_fd_sc_hd__xor2_2 _19263_ (.A(_14285_),
    .B(_14428_),
    .X(_14439_));
 sky130_fd_sc_hd__nand2_2 _19264_ (.A(_13683_),
    .B(_13793_),
    .Y(_14450_));
 sky130_fd_sc_hd__xnor2_2 _19265_ (.A(_14439_),
    .B(_14450_),
    .Y(_14461_));
 sky130_fd_sc_hd__xnor2_2 _19266_ (.A(_13760_),
    .B(_14461_),
    .Y(_14472_));
 sky130_fd_sc_hd__a21bo_2 _19267_ (.A1(_13180_),
    .A2(_13826_),
    .B1_N(_13815_),
    .X(_14483_));
 sky130_fd_sc_hd__xnor2_2 _19268_ (.A(_14472_),
    .B(_14483_),
    .Y(_14494_));
 sky130_fd_sc_hd__nor3_2 _19269_ (.A(_13235_),
    .B(_13837_),
    .C(_13848_),
    .Y(_14505_));
 sky130_fd_sc_hd__a21oi_2 _19270_ (.A1(_13257_),
    .A2(_13870_),
    .B1(_14505_),
    .Y(_14515_));
 sky130_fd_sc_hd__xnor2_2 _19271_ (.A(_14494_),
    .B(_14515_),
    .Y(_14526_));
 sky130_fd_sc_hd__nor3_2 _19272_ (.A(_13978_),
    .B(_13989_),
    .C(_14526_),
    .Y(_14537_));
 sky130_fd_sc_hd__o21a_2 _19273_ (.A1(_13978_),
    .A2(_13989_),
    .B1(_14526_),
    .X(_14548_));
 sky130_fd_sc_hd__nor2_2 _19274_ (.A(_14537_),
    .B(_14548_),
    .Y(_14559_));
 sky130_fd_sc_hd__o21ba_2 _19275_ (.A1(_13935_),
    .A2(_13957_),
    .B1_N(_13924_),
    .X(_14570_));
 sky130_fd_sc_hd__xnor2_2 _19276_ (.A(_14559_),
    .B(_14570_),
    .Y(oO[11]));
 sky130_fd_sc_hd__nor2_2 _19277_ (.A(_13859_),
    .B(_14494_),
    .Y(_14591_));
 sky130_fd_sc_hd__nand2_2 _19278_ (.A(_14472_),
    .B(_14483_),
    .Y(_14602_));
 sky130_fd_sc_hd__nand2_2 _19279_ (.A(_14439_),
    .B(_14450_),
    .Y(_14613_));
 sky130_fd_sc_hd__nand2_2 _19280_ (.A(_13705_),
    .B(_13716_),
    .Y(_14624_));
 sky130_fd_sc_hd__or3b_2 _19281_ (.A(_13749_),
    .B(_14461_),
    .C_N(_14624_),
    .X(_14635_));
 sky130_fd_sc_hd__or2b_2 _19282_ (.A(_14263_),
    .B_N(_14274_),
    .X(_14646_));
 sky130_fd_sc_hd__nand2_2 _19283_ (.A(_14285_),
    .B(_14428_),
    .Y(_14657_));
 sky130_fd_sc_hd__or2_2 _19284_ (.A(_14132_),
    .B(_14143_),
    .X(_14668_));
 sky130_fd_sc_hd__nand2_2 _19285_ (.A(_14154_),
    .B(_14252_),
    .Y(_14679_));
 sky130_fd_sc_hd__nand2_2 _19286_ (.A(_14044_),
    .B(_14055_),
    .Y(_14690_));
 sky130_fd_sc_hd__nand2_2 _19287_ (.A(_14066_),
    .B(_14121_),
    .Y(_14701_));
 sky130_fd_sc_hd__and4_2 _19288_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[11]),
    .D(iX[12]),
    .X(_14712_));
 sky130_fd_sc_hd__a22oi_2 _19289_ (.A1(iY[1]),
    .A2(iX[11]),
    .B1(iX[12]),
    .B2(iY[0]),
    .Y(_14723_));
 sky130_fd_sc_hd__nor2_2 _19290_ (.A(_14712_),
    .B(_14723_),
    .Y(_14734_));
 sky130_fd_sc_hd__nand2_2 _19291_ (.A(iY[2]),
    .B(iX[10]),
    .Y(_14745_));
 sky130_fd_sc_hd__xnor2_2 _19292_ (.A(_14734_),
    .B(_14745_),
    .Y(_14756_));
 sky130_fd_sc_hd__o21ba_2 _19293_ (.A1(_14011_),
    .A2(_14033_),
    .B1_N(_14000_),
    .X(_14767_));
 sky130_fd_sc_hd__xnor2_2 _19294_ (.A(_14756_),
    .B(_14767_),
    .Y(_14778_));
 sky130_fd_sc_hd__and4_2 _19295_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[8]),
    .D(iX[9]),
    .X(_14789_));
 sky130_fd_sc_hd__a22oi_2 _19296_ (.A1(iY[4]),
    .A2(iX[8]),
    .B1(iX[9]),
    .B2(iY[3]),
    .Y(_14800_));
 sky130_fd_sc_hd__nor2_2 _19297_ (.A(_14789_),
    .B(_14800_),
    .Y(_14811_));
 sky130_fd_sc_hd__nand2_2 _19298_ (.A(iY[5]),
    .B(iX[7]),
    .Y(_14822_));
 sky130_fd_sc_hd__xnor2_2 _19299_ (.A(_14811_),
    .B(_14822_),
    .Y(_14832_));
 sky130_fd_sc_hd__xnor2_2 _19300_ (.A(_14778_),
    .B(_14832_),
    .Y(_14843_));
 sky130_fd_sc_hd__a21o_2 _19301_ (.A1(_14690_),
    .A2(_14701_),
    .B1(_14843_),
    .X(_14854_));
 sky130_fd_sc_hd__nand3_2 _19302_ (.A(_14690_),
    .B(_14701_),
    .C(_14843_),
    .Y(_14865_));
 sky130_fd_sc_hd__o21ba_2 _19303_ (.A1(_14198_),
    .A2(_14219_),
    .B1_N(_14187_),
    .X(_14876_));
 sky130_fd_sc_hd__o21ba_2 _19304_ (.A1(_14088_),
    .A2(_14110_),
    .B1_N(_14077_),
    .X(_14887_));
 sky130_fd_sc_hd__and4_2 _19305_ (.A(iX[5]),
    .B(iX[6]),
    .C(iY[6]),
    .D(iY[7]),
    .X(_14898_));
 sky130_fd_sc_hd__a22oi_2 _19306_ (.A1(iX[6]),
    .A2(iY[6]),
    .B1(iY[7]),
    .B2(iX[5]),
    .Y(_14909_));
 sky130_fd_sc_hd__nor2_2 _19307_ (.A(_14898_),
    .B(_14909_),
    .Y(_14920_));
 sky130_fd_sc_hd__nand2_2 _19308_ (.A(iX[4]),
    .B(iY[8]),
    .Y(_14931_));
 sky130_fd_sc_hd__xnor2_2 _19309_ (.A(_14920_),
    .B(_14931_),
    .Y(_14942_));
 sky130_fd_sc_hd__xnor2_2 _19310_ (.A(_14887_),
    .B(_14942_),
    .Y(_14953_));
 sky130_fd_sc_hd__xnor2_2 _19311_ (.A(_14876_),
    .B(_14953_),
    .Y(_14964_));
 sky130_fd_sc_hd__and3_2 _19312_ (.A(_14854_),
    .B(_14865_),
    .C(_14964_),
    .X(_14975_));
 sky130_fd_sc_hd__a21oi_2 _19313_ (.A1(_14854_),
    .A2(_14865_),
    .B1(_14964_),
    .Y(_14986_));
 sky130_fd_sc_hd__a211oi_2 _19314_ (.A1(_14668_),
    .A2(_14679_),
    .B1(_14975_),
    .C1(_14986_),
    .Y(_14997_));
 sky130_fd_sc_hd__o211a_2 _19315_ (.A1(_14975_),
    .A2(_14986_),
    .B1(_14668_),
    .C1(_14679_),
    .X(_15008_));
 sky130_fd_sc_hd__or2b_2 _19316_ (.A(_14176_),
    .B_N(_14230_),
    .X(_15019_));
 sky130_fd_sc_hd__or2b_2 _19317_ (.A(_14165_),
    .B_N(_14241_),
    .X(_15030_));
 sky130_fd_sc_hd__nand2_2 _19318_ (.A(_15019_),
    .B(_15030_),
    .Y(_15041_));
 sky130_fd_sc_hd__and4_2 _19319_ (.A(iX[2]),
    .B(iX[3]),
    .C(iY[9]),
    .D(iY[10]),
    .X(_15052_));
 sky130_fd_sc_hd__a22oi_2 _19320_ (.A1(iX[3]),
    .A2(iY[9]),
    .B1(iY[10]),
    .B2(iX[2]),
    .Y(_15063_));
 sky130_fd_sc_hd__nor2_2 _19321_ (.A(_15052_),
    .B(_15063_),
    .Y(_15074_));
 sky130_fd_sc_hd__nand2_2 _19322_ (.A(iX[1]),
    .B(iY[11]),
    .Y(_15085_));
 sky130_fd_sc_hd__xnor2_2 _19323_ (.A(_15074_),
    .B(_15085_),
    .Y(_15096_));
 sky130_fd_sc_hd__o21ba_2 _19324_ (.A1(_14329_),
    .A2(_14351_),
    .B1_N(_14318_),
    .X(_15107_));
 sky130_fd_sc_hd__xnor2_2 _19325_ (.A(_15096_),
    .B(_15107_),
    .Y(_15118_));
 sky130_fd_sc_hd__and2_2 _19326_ (.A(iX[0]),
    .B(iY[12]),
    .X(_15129_));
 sky130_fd_sc_hd__nor2_2 _19327_ (.A(_15118_),
    .B(_15129_),
    .Y(_15139_));
 sky130_fd_sc_hd__and2_2 _19328_ (.A(_15118_),
    .B(_15129_),
    .X(_15150_));
 sky130_fd_sc_hd__or2_2 _19329_ (.A(_15139_),
    .B(_15150_),
    .X(_15161_));
 sky130_fd_sc_hd__xnor2_2 _19330_ (.A(_15041_),
    .B(_15161_),
    .Y(_15172_));
 sky130_fd_sc_hd__xnor2_2 _19331_ (.A(_14373_),
    .B(_15172_),
    .Y(_15183_));
 sky130_fd_sc_hd__o21a_2 _19332_ (.A1(_14997_),
    .A2(_15008_),
    .B1(_15183_),
    .X(_15194_));
 sky130_fd_sc_hd__nor3_2 _19333_ (.A(_14997_),
    .B(_15008_),
    .C(_15183_),
    .Y(_15205_));
 sky130_fd_sc_hd__a211oi_2 _19334_ (.A1(_14646_),
    .A2(_14657_),
    .B1(_15194_),
    .C1(_15205_),
    .Y(_15216_));
 sky130_fd_sc_hd__o211a_2 _19335_ (.A1(_15194_),
    .A2(_15205_),
    .B1(_14646_),
    .C1(_14657_),
    .X(_15227_));
 sky130_fd_sc_hd__o21ba_2 _19336_ (.A1(_15216_),
    .A2(_15227_),
    .B1_N(_14406_),
    .X(_15238_));
 sky130_fd_sc_hd__nor3b_2 _19337_ (.A(_15216_),
    .B(_15227_),
    .C_N(_14406_),
    .Y(_15249_));
 sky130_fd_sc_hd__a211oi_2 _19338_ (.A1(_14613_),
    .A2(_14635_),
    .B1(_15238_),
    .C1(_15249_),
    .Y(_15260_));
 sky130_fd_sc_hd__o211a_2 _19339_ (.A1(_15238_),
    .A2(_15249_),
    .B1(_14613_),
    .C1(_14635_),
    .X(_15271_));
 sky130_fd_sc_hd__or3_2 _19340_ (.A(_14602_),
    .B(_15260_),
    .C(_15271_),
    .X(_15282_));
 sky130_fd_sc_hd__o21ai_2 _19341_ (.A1(_15260_),
    .A2(_15271_),
    .B1(_14602_),
    .Y(_15293_));
 sky130_fd_sc_hd__and3_2 _19342_ (.A(_14591_),
    .B(_15282_),
    .C(_15293_),
    .X(_15304_));
 sky130_fd_sc_hd__a21oi_2 _19343_ (.A1(_15282_),
    .A2(_15293_),
    .B1(_14591_),
    .Y(_15315_));
 sky130_fd_sc_hd__and4bb_2 _19344_ (.A_N(_14505_),
    .B_N(_14494_),
    .C(_13870_),
    .D(_13257_),
    .X(_15326_));
 sky130_fd_sc_hd__nor3b_2 _19345_ (.A(_15304_),
    .B(_15315_),
    .C_N(_15326_),
    .Y(_15337_));
 sky130_fd_sc_hd__o21bai_2 _19346_ (.A1(_15304_),
    .A2(_15315_),
    .B1_N(_15326_),
    .Y(_15348_));
 sky130_fd_sc_hd__or2b_2 _19347_ (.A(_15337_),
    .B_N(_15348_),
    .X(_15359_));
 sky130_fd_sc_hd__o21bai_2 _19348_ (.A1(_14548_),
    .A2(_14570_),
    .B1_N(_14537_),
    .Y(_15370_));
 sky130_fd_sc_hd__xnor2_2 _19349_ (.A(_15359_),
    .B(_15370_),
    .Y(oO[12]));
 sky130_fd_sc_hd__a21o_2 _19350_ (.A1(_15348_),
    .A2(_15370_),
    .B1(_15337_),
    .X(_15391_));
 sky130_fd_sc_hd__nand3_2 _19351_ (.A(_14854_),
    .B(_14865_),
    .C(_14964_),
    .Y(_15402_));
 sky130_fd_sc_hd__or2b_2 _19352_ (.A(_14767_),
    .B_N(_14756_),
    .X(_15413_));
 sky130_fd_sc_hd__nand2_2 _19353_ (.A(_14778_),
    .B(_14832_),
    .Y(_15424_));
 sky130_fd_sc_hd__and4_2 _19354_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[12]),
    .D(iX[13]),
    .X(_15435_));
 sky130_fd_sc_hd__a22oi_2 _19355_ (.A1(iY[1]),
    .A2(iX[12]),
    .B1(iX[13]),
    .B2(iY[0]),
    .Y(_15446_));
 sky130_fd_sc_hd__nor2_2 _19356_ (.A(_15435_),
    .B(_15446_),
    .Y(_15457_));
 sky130_fd_sc_hd__nand2_2 _19357_ (.A(iY[2]),
    .B(iX[11]),
    .Y(_15467_));
 sky130_fd_sc_hd__xnor2_2 _19358_ (.A(_15457_),
    .B(_15467_),
    .Y(_15478_));
 sky130_fd_sc_hd__o21ba_2 _19359_ (.A1(_14723_),
    .A2(_14745_),
    .B1_N(_14712_),
    .X(_15489_));
 sky130_fd_sc_hd__xnor2_2 _19360_ (.A(_15478_),
    .B(_15489_),
    .Y(_15500_));
 sky130_fd_sc_hd__and4_2 _19361_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[9]),
    .D(iX[10]),
    .X(_15511_));
 sky130_fd_sc_hd__a22oi_2 _19362_ (.A1(iY[4]),
    .A2(iX[9]),
    .B1(iX[10]),
    .B2(iY[3]),
    .Y(_15522_));
 sky130_fd_sc_hd__nor2_2 _19363_ (.A(_15511_),
    .B(_15522_),
    .Y(_15533_));
 sky130_fd_sc_hd__nand2_2 _19364_ (.A(iY[5]),
    .B(iX[8]),
    .Y(_15544_));
 sky130_fd_sc_hd__xnor2_2 _19365_ (.A(_15533_),
    .B(_15544_),
    .Y(_15555_));
 sky130_fd_sc_hd__xnor2_2 _19366_ (.A(_15500_),
    .B(_15555_),
    .Y(_15566_));
 sky130_fd_sc_hd__a21o_2 _19367_ (.A1(_15413_),
    .A2(_15424_),
    .B1(_15566_),
    .X(_15577_));
 sky130_fd_sc_hd__nand3_2 _19368_ (.A(_15413_),
    .B(_15424_),
    .C(_15566_),
    .Y(_15588_));
 sky130_fd_sc_hd__o21ba_2 _19369_ (.A1(_14909_),
    .A2(_14931_),
    .B1_N(_14898_),
    .X(_15599_));
 sky130_fd_sc_hd__o21ba_2 _19370_ (.A1(_14800_),
    .A2(_14822_),
    .B1_N(_14789_),
    .X(_15610_));
 sky130_fd_sc_hd__and4_2 _19371_ (.A(iX[6]),
    .B(iY[6]),
    .C(iX[7]),
    .D(iY[7]),
    .X(_15621_));
 sky130_fd_sc_hd__a22oi_2 _19372_ (.A1(iY[6]),
    .A2(iX[7]),
    .B1(iY[7]),
    .B2(iX[6]),
    .Y(_15632_));
 sky130_fd_sc_hd__nor2_2 _19373_ (.A(_15621_),
    .B(_15632_),
    .Y(_15643_));
 sky130_fd_sc_hd__nand2_2 _19374_ (.A(iX[5]),
    .B(iY[8]),
    .Y(_15654_));
 sky130_fd_sc_hd__xnor2_2 _19375_ (.A(_15643_),
    .B(_15654_),
    .Y(_15665_));
 sky130_fd_sc_hd__xnor2_2 _19376_ (.A(_15610_),
    .B(_15665_),
    .Y(_15676_));
 sky130_fd_sc_hd__xnor2_2 _19377_ (.A(_15599_),
    .B(_15676_),
    .Y(_15687_));
 sky130_fd_sc_hd__and3_2 _19378_ (.A(_15577_),
    .B(_15588_),
    .C(_15687_),
    .X(_15698_));
 sky130_fd_sc_hd__a21oi_2 _19379_ (.A1(_15577_),
    .A2(_15588_),
    .B1(_15687_),
    .Y(_15709_));
 sky130_fd_sc_hd__a211o_2 _19380_ (.A1(_14854_),
    .A2(_15402_),
    .B1(_15698_),
    .C1(_15709_),
    .X(_15720_));
 sky130_fd_sc_hd__o211ai_2 _19381_ (.A1(_15698_),
    .A2(_15709_),
    .B1(_14854_),
    .C1(_15402_),
    .Y(_15731_));
 sky130_fd_sc_hd__and2b_2 _19382_ (.A_N(_15107_),
    .B(_15096_),
    .X(_15742_));
 sky130_fd_sc_hd__and2b_2 _19383_ (.A_N(_14887_),
    .B(_14942_),
    .X(_15753_));
 sky130_fd_sc_hd__and2b_2 _19384_ (.A_N(_14876_),
    .B(_14953_),
    .X(_15764_));
 sky130_fd_sc_hd__a22oi_2 _19385_ (.A1(iX[1]),
    .A2(iY[12]),
    .B1(iY[13]),
    .B2(iX[0]),
    .Y(_15775_));
 sky130_fd_sc_hd__and3_2 _19386_ (.A(iX[1]),
    .B(iY[13]),
    .C(_15129_),
    .X(_15786_));
 sky130_fd_sc_hd__or2_2 _19387_ (.A(_15775_),
    .B(_15786_),
    .X(_15797_));
 sky130_fd_sc_hd__and4_2 _19388_ (.A(iX[3]),
    .B(iX[4]),
    .C(iY[9]),
    .D(iY[10]),
    .X(_15808_));
 sky130_fd_sc_hd__a22oi_2 _19389_ (.A1(iX[4]),
    .A2(iY[9]),
    .B1(iY[10]),
    .B2(iX[3]),
    .Y(_15819_));
 sky130_fd_sc_hd__nor2_2 _19390_ (.A(_15808_),
    .B(_15819_),
    .Y(_15829_));
 sky130_fd_sc_hd__nand2_2 _19391_ (.A(iX[2]),
    .B(iY[11]),
    .Y(_15840_));
 sky130_fd_sc_hd__xnor2_2 _19392_ (.A(_15829_),
    .B(_15840_),
    .Y(_15851_));
 sky130_fd_sc_hd__o21ba_2 _19393_ (.A1(_15063_),
    .A2(_15085_),
    .B1_N(_15052_),
    .X(_15862_));
 sky130_fd_sc_hd__xnor2_2 _19394_ (.A(_15851_),
    .B(_15862_),
    .Y(_15873_));
 sky130_fd_sc_hd__xnor2_2 _19395_ (.A(_15797_),
    .B(_15873_),
    .Y(_15884_));
 sky130_fd_sc_hd__o21ai_2 _19396_ (.A1(_15753_),
    .A2(_15764_),
    .B1(_15884_),
    .Y(_15895_));
 sky130_fd_sc_hd__or3_2 _19397_ (.A(_15753_),
    .B(_15764_),
    .C(_15884_),
    .X(_15906_));
 sky130_fd_sc_hd__o211a_2 _19398_ (.A1(_15742_),
    .A2(_15150_),
    .B1(_15895_),
    .C1(_15906_),
    .X(_15917_));
 sky130_fd_sc_hd__inv_2 _19399_ (.A(_15917_),
    .Y(_15928_));
 sky130_fd_sc_hd__a211o_2 _19400_ (.A1(_15895_),
    .A2(_15906_),
    .B1(_15742_),
    .C1(_15150_),
    .X(_15939_));
 sky130_fd_sc_hd__nand4_2 _19401_ (.A(_15720_),
    .B(_15731_),
    .C(_15928_),
    .D(_15939_),
    .Y(_15950_));
 sky130_fd_sc_hd__a22o_2 _19402_ (.A1(_15720_),
    .A2(_15731_),
    .B1(_15928_),
    .B2(_15939_),
    .X(_15961_));
 sky130_fd_sc_hd__nand2_2 _19403_ (.A(_15950_),
    .B(_15961_),
    .Y(_15972_));
 sky130_fd_sc_hd__or2_2 _19404_ (.A(_14997_),
    .B(_15205_),
    .X(_15983_));
 sky130_fd_sc_hd__xor2_2 _19405_ (.A(_15972_),
    .B(_15983_),
    .X(_15994_));
 sky130_fd_sc_hd__and2b_2 _19406_ (.A_N(_15161_),
    .B(_15041_),
    .X(_16005_));
 sky130_fd_sc_hd__a21oi_2 _19407_ (.A1(_14373_),
    .A2(_15172_),
    .B1(_16005_),
    .Y(_16016_));
 sky130_fd_sc_hd__xnor2_2 _19408_ (.A(_15994_),
    .B(_16016_),
    .Y(_16027_));
 sky130_fd_sc_hd__or2_2 _19409_ (.A(_15216_),
    .B(_15249_),
    .X(_16038_));
 sky130_fd_sc_hd__xnor2_2 _19410_ (.A(_16027_),
    .B(_16038_),
    .Y(_16049_));
 sky130_fd_sc_hd__xnor2_2 _19411_ (.A(_15260_),
    .B(_16049_),
    .Y(_16060_));
 sky130_fd_sc_hd__a21bo_2 _19412_ (.A1(_14591_),
    .A2(_15293_),
    .B1_N(_15282_),
    .X(_16071_));
 sky130_fd_sc_hd__xnor2_2 _19413_ (.A(_16060_),
    .B(_16071_),
    .Y(_16082_));
 sky130_fd_sc_hd__xor2_2 _19414_ (.A(_15391_),
    .B(_16082_),
    .X(oO[13]));
 sky130_fd_sc_hd__inv_2 _19415_ (.A(_15304_),
    .Y(_16103_));
 sky130_fd_sc_hd__a2bb2o_2 _19416_ (.A1_N(_16103_),
    .A2_N(_16060_),
    .B1(_16082_),
    .B2(_15391_),
    .X(_16114_));
 sky130_fd_sc_hd__and2b_2 _19417_ (.A_N(_16027_),
    .B(_16038_),
    .X(_16125_));
 sky130_fd_sc_hd__nand3_2 _19418_ (.A(_15577_),
    .B(_15588_),
    .C(_15687_),
    .Y(_16136_));
 sky130_fd_sc_hd__or2b_2 _19419_ (.A(_15489_),
    .B_N(_15478_),
    .X(_16146_));
 sky130_fd_sc_hd__nand2_2 _19420_ (.A(_15500_),
    .B(_15555_),
    .Y(_16157_));
 sky130_fd_sc_hd__and4_2 _19421_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[13]),
    .D(iX[14]),
    .X(_16168_));
 sky130_fd_sc_hd__a22oi_2 _19422_ (.A1(iY[1]),
    .A2(iX[13]),
    .B1(iX[14]),
    .B2(iY[0]),
    .Y(_16179_));
 sky130_fd_sc_hd__nor2_2 _19423_ (.A(_16168_),
    .B(_16179_),
    .Y(_16190_));
 sky130_fd_sc_hd__nand2_2 _19424_ (.A(iY[2]),
    .B(iX[12]),
    .Y(_16201_));
 sky130_fd_sc_hd__xnor2_2 _19425_ (.A(_16190_),
    .B(_16201_),
    .Y(_16212_));
 sky130_fd_sc_hd__o21ba_2 _19426_ (.A1(_15446_),
    .A2(_15467_),
    .B1_N(_15435_),
    .X(_16223_));
 sky130_fd_sc_hd__xnor2_2 _19427_ (.A(_16212_),
    .B(_16223_),
    .Y(_16234_));
 sky130_fd_sc_hd__and4_2 _19428_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[10]),
    .D(iX[11]),
    .X(_16245_));
 sky130_fd_sc_hd__a22oi_2 _19429_ (.A1(iY[4]),
    .A2(iX[10]),
    .B1(iX[11]),
    .B2(iY[3]),
    .Y(_16256_));
 sky130_fd_sc_hd__nor2_2 _19430_ (.A(_16245_),
    .B(_16256_),
    .Y(_16267_));
 sky130_fd_sc_hd__nand2_2 _19431_ (.A(iY[5]),
    .B(iX[9]),
    .Y(_16278_));
 sky130_fd_sc_hd__xnor2_2 _19432_ (.A(_16267_),
    .B(_16278_),
    .Y(_16289_));
 sky130_fd_sc_hd__xnor2_2 _19433_ (.A(_16234_),
    .B(_16289_),
    .Y(_16300_));
 sky130_fd_sc_hd__a21o_2 _19434_ (.A1(_16146_),
    .A2(_16157_),
    .B1(_16300_),
    .X(_16311_));
 sky130_fd_sc_hd__nand3_2 _19435_ (.A(_16146_),
    .B(_16157_),
    .C(_16300_),
    .Y(_16322_));
 sky130_fd_sc_hd__o21ba_2 _19436_ (.A1(_15632_),
    .A2(_15654_),
    .B1_N(_15621_),
    .X(_16333_));
 sky130_fd_sc_hd__o21ba_2 _19437_ (.A1(_15522_),
    .A2(_15544_),
    .B1_N(_15511_),
    .X(_16344_));
 sky130_fd_sc_hd__and4_2 _19438_ (.A(iY[6]),
    .B(iX[7]),
    .C(iY[7]),
    .D(iX[8]),
    .X(_16355_));
 sky130_fd_sc_hd__a22oi_2 _19439_ (.A1(iX[7]),
    .A2(iY[7]),
    .B1(iX[8]),
    .B2(iY[6]),
    .Y(_16366_));
 sky130_fd_sc_hd__nor2_2 _19440_ (.A(_16355_),
    .B(_16366_),
    .Y(_16377_));
 sky130_fd_sc_hd__nand2_2 _19441_ (.A(iX[6]),
    .B(iY[8]),
    .Y(_16388_));
 sky130_fd_sc_hd__xnor2_2 _19442_ (.A(_16377_),
    .B(_16388_),
    .Y(_16399_));
 sky130_fd_sc_hd__xnor2_2 _19443_ (.A(_16344_),
    .B(_16399_),
    .Y(_16410_));
 sky130_fd_sc_hd__xnor2_2 _19444_ (.A(_16333_),
    .B(_16410_),
    .Y(_16421_));
 sky130_fd_sc_hd__nand3_2 _19445_ (.A(_16311_),
    .B(_16322_),
    .C(_16421_),
    .Y(_16432_));
 sky130_fd_sc_hd__a21o_2 _19446_ (.A1(_16311_),
    .A2(_16322_),
    .B1(_16421_),
    .X(_16443_));
 sky130_fd_sc_hd__nand2_2 _19447_ (.A(_16432_),
    .B(_16443_),
    .Y(_16454_));
 sky130_fd_sc_hd__a21o_2 _19448_ (.A1(_15577_),
    .A2(_16136_),
    .B1(_16454_),
    .X(_16465_));
 sky130_fd_sc_hd__nand3_2 _19449_ (.A(_15577_),
    .B(_16136_),
    .C(_16454_),
    .Y(_16476_));
 sky130_fd_sc_hd__or2b_2 _19450_ (.A(_15862_),
    .B_N(_15851_),
    .X(_16486_));
 sky130_fd_sc_hd__or2b_2 _19451_ (.A(_15797_),
    .B_N(_15873_),
    .X(_16497_));
 sky130_fd_sc_hd__or2b_2 _19452_ (.A(_15610_),
    .B_N(_15665_),
    .X(_16508_));
 sky130_fd_sc_hd__or2b_2 _19453_ (.A(_15599_),
    .B_N(_15676_),
    .X(_16519_));
 sky130_fd_sc_hd__and4_2 _19454_ (.A(iX[1]),
    .B(iX[2]),
    .C(iY[12]),
    .D(iY[13]),
    .X(_16530_));
 sky130_fd_sc_hd__a22oi_2 _19455_ (.A1(iX[2]),
    .A2(iY[12]),
    .B1(iY[13]),
    .B2(iX[1]),
    .Y(_16541_));
 sky130_fd_sc_hd__nor2_2 _19456_ (.A(_16530_),
    .B(_16541_),
    .Y(_16552_));
 sky130_fd_sc_hd__nand2_2 _19457_ (.A(iX[0]),
    .B(iY[14]),
    .Y(_16563_));
 sky130_fd_sc_hd__xnor2_2 _19458_ (.A(_16552_),
    .B(_16563_),
    .Y(_16574_));
 sky130_fd_sc_hd__and4_2 _19459_ (.A(iX[4]),
    .B(iX[5]),
    .C(iY[9]),
    .D(iY[10]),
    .X(_16585_));
 sky130_fd_sc_hd__a22oi_2 _19460_ (.A1(iX[5]),
    .A2(iY[9]),
    .B1(iY[10]),
    .B2(iX[4]),
    .Y(_16596_));
 sky130_fd_sc_hd__nor2_2 _19461_ (.A(_16585_),
    .B(_16596_),
    .Y(_16607_));
 sky130_fd_sc_hd__nand2_2 _19462_ (.A(iX[3]),
    .B(iY[11]),
    .Y(_16618_));
 sky130_fd_sc_hd__xnor2_2 _19463_ (.A(_16607_),
    .B(_16618_),
    .Y(_16629_));
 sky130_fd_sc_hd__o21ba_2 _19464_ (.A1(_15819_),
    .A2(_15840_),
    .B1_N(_15808_),
    .X(_16640_));
 sky130_fd_sc_hd__xnor2_2 _19465_ (.A(_16629_),
    .B(_16640_),
    .Y(_16651_));
 sky130_fd_sc_hd__and2_2 _19466_ (.A(_16574_),
    .B(_16651_),
    .X(_16662_));
 sky130_fd_sc_hd__nor2_2 _19467_ (.A(_16574_),
    .B(_16651_),
    .Y(_16673_));
 sky130_fd_sc_hd__or2_2 _19468_ (.A(_16662_),
    .B(_16673_),
    .X(_16684_));
 sky130_fd_sc_hd__a21o_2 _19469_ (.A1(_16508_),
    .A2(_16519_),
    .B1(_16684_),
    .X(_16695_));
 sky130_fd_sc_hd__inv_2 _19470_ (.A(_16695_),
    .Y(_16706_));
 sky130_fd_sc_hd__and3_2 _19471_ (.A(_16508_),
    .B(_16519_),
    .C(_16684_),
    .X(_16717_));
 sky130_fd_sc_hd__a211o_2 _19472_ (.A1(_16486_),
    .A2(_16497_),
    .B1(_16706_),
    .C1(_16717_),
    .X(_16728_));
 sky130_fd_sc_hd__o211ai_2 _19473_ (.A1(_16706_),
    .A2(_16717_),
    .B1(_16486_),
    .C1(_16497_),
    .Y(_16739_));
 sky130_fd_sc_hd__and4_2 _19474_ (.A(_16465_),
    .B(_16476_),
    .C(_16728_),
    .D(_16739_),
    .X(_16750_));
 sky130_fd_sc_hd__a22oi_2 _19475_ (.A1(_16465_),
    .A2(_16476_),
    .B1(_16728_),
    .B2(_16739_),
    .Y(_16761_));
 sky130_fd_sc_hd__a211o_2 _19476_ (.A1(_15720_),
    .A2(_15950_),
    .B1(_16750_),
    .C1(_16761_),
    .X(_16772_));
 sky130_fd_sc_hd__o211ai_2 _19477_ (.A1(_16750_),
    .A2(_16761_),
    .B1(_15720_),
    .C1(_15950_),
    .Y(_16783_));
 sky130_fd_sc_hd__o21a_2 _19478_ (.A1(_15753_),
    .A2(_15764_),
    .B1(_15884_),
    .X(_16794_));
 sky130_fd_sc_hd__o21ai_2 _19479_ (.A1(_16794_),
    .A2(_15917_),
    .B1(_15786_),
    .Y(_16805_));
 sky130_fd_sc_hd__or3_2 _19480_ (.A(_15786_),
    .B(_16794_),
    .C(_15917_),
    .X(_16815_));
 sky130_fd_sc_hd__and2_2 _19481_ (.A(_16805_),
    .B(_16815_),
    .X(_16826_));
 sky130_fd_sc_hd__a21oi_2 _19482_ (.A1(_16772_),
    .A2(_16783_),
    .B1(_16826_),
    .Y(_16837_));
 sky130_fd_sc_hd__and3_2 _19483_ (.A(_16772_),
    .B(_16783_),
    .C(_16826_),
    .X(_16848_));
 sky130_fd_sc_hd__nor2_2 _19484_ (.A(_16837_),
    .B(_16848_),
    .Y(_16859_));
 sky130_fd_sc_hd__or2b_2 _19485_ (.A(_15972_),
    .B_N(_15983_),
    .X(_16870_));
 sky130_fd_sc_hd__o21a_2 _19486_ (.A1(_15994_),
    .A2(_16016_),
    .B1(_16870_),
    .X(_16881_));
 sky130_fd_sc_hd__xor2_2 _19487_ (.A(_16859_),
    .B(_16881_),
    .X(_16892_));
 sky130_fd_sc_hd__xor2_2 _19488_ (.A(_16125_),
    .B(_16892_),
    .X(_16903_));
 sky130_fd_sc_hd__nand2_2 _19489_ (.A(_15260_),
    .B(_16049_),
    .Y(_16914_));
 sky130_fd_sc_hd__or2_2 _19490_ (.A(_15282_),
    .B(_16060_),
    .X(_16925_));
 sky130_fd_sc_hd__nand2_2 _19491_ (.A(_16914_),
    .B(_16925_),
    .Y(_16936_));
 sky130_fd_sc_hd__xnor2_2 _19492_ (.A(_16903_),
    .B(_16936_),
    .Y(_16947_));
 sky130_fd_sc_hd__xor2_2 _19493_ (.A(_16114_),
    .B(_16947_),
    .X(oO[14]));
 sky130_fd_sc_hd__a2bb2o_2 _19494_ (.A1_N(_16925_),
    .A2_N(_16903_),
    .B1(_16947_),
    .B2(_16114_),
    .X(_16968_));
 sky130_fd_sc_hd__or3_2 _19495_ (.A(_16837_),
    .B(_16848_),
    .C(_16881_),
    .X(_16979_));
 sky130_fd_sc_hd__inv_2 _19496_ (.A(_16465_),
    .Y(_16990_));
 sky130_fd_sc_hd__or2b_2 _19497_ (.A(_16223_),
    .B_N(_16212_),
    .X(_17001_));
 sky130_fd_sc_hd__nand2_2 _19498_ (.A(_16234_),
    .B(_16289_),
    .Y(_17012_));
 sky130_fd_sc_hd__and4_2 _19499_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[14]),
    .D(iX[15]),
    .X(_17023_));
 sky130_fd_sc_hd__a22oi_2 _19500_ (.A1(iY[1]),
    .A2(iX[14]),
    .B1(iX[15]),
    .B2(iY[0]),
    .Y(_17034_));
 sky130_fd_sc_hd__nor2_2 _19501_ (.A(_17023_),
    .B(_17034_),
    .Y(_17045_));
 sky130_fd_sc_hd__nand2_2 _19502_ (.A(iY[2]),
    .B(iX[13]),
    .Y(_17056_));
 sky130_fd_sc_hd__xnor2_2 _19503_ (.A(_17045_),
    .B(_17056_),
    .Y(_17067_));
 sky130_fd_sc_hd__o21ba_2 _19504_ (.A1(_16179_),
    .A2(_16201_),
    .B1_N(_16168_),
    .X(_17078_));
 sky130_fd_sc_hd__xnor2_2 _19505_ (.A(_17067_),
    .B(_17078_),
    .Y(_17089_));
 sky130_fd_sc_hd__and4_2 _19506_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[11]),
    .D(iX[12]),
    .X(_17100_));
 sky130_fd_sc_hd__a22oi_2 _19507_ (.A1(iY[4]),
    .A2(iX[11]),
    .B1(iX[12]),
    .B2(iY[3]),
    .Y(_17111_));
 sky130_fd_sc_hd__nor2_2 _19508_ (.A(_17100_),
    .B(_17111_),
    .Y(_17122_));
 sky130_fd_sc_hd__nand2_2 _19509_ (.A(iY[5]),
    .B(iX[10]),
    .Y(_17133_));
 sky130_fd_sc_hd__xnor2_2 _19510_ (.A(_17122_),
    .B(_17133_),
    .Y(_17144_));
 sky130_fd_sc_hd__xnor2_2 _19511_ (.A(_17089_),
    .B(_17144_),
    .Y(_17155_));
 sky130_fd_sc_hd__a21o_2 _19512_ (.A1(_17001_),
    .A2(_17012_),
    .B1(_17155_),
    .X(_17166_));
 sky130_fd_sc_hd__nand3_2 _19513_ (.A(_17001_),
    .B(_17012_),
    .C(_17155_),
    .Y(_17177_));
 sky130_fd_sc_hd__o21ba_2 _19514_ (.A1(_16366_),
    .A2(_16388_),
    .B1_N(_16355_),
    .X(_17188_));
 sky130_fd_sc_hd__o21ba_2 _19515_ (.A1(_16256_),
    .A2(_16278_),
    .B1_N(_16245_),
    .X(_17198_));
 sky130_fd_sc_hd__and4_2 _19516_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[8]),
    .D(iX[9]),
    .X(_17209_));
 sky130_fd_sc_hd__a22oi_2 _19517_ (.A1(iY[7]),
    .A2(iX[8]),
    .B1(iX[9]),
    .B2(iY[6]),
    .Y(_17220_));
 sky130_fd_sc_hd__nor2_2 _19518_ (.A(_17209_),
    .B(_17220_),
    .Y(_17231_));
 sky130_fd_sc_hd__nand2_2 _19519_ (.A(iX[7]),
    .B(iY[8]),
    .Y(_17242_));
 sky130_fd_sc_hd__xnor2_2 _19520_ (.A(_17231_),
    .B(_17242_),
    .Y(_17253_));
 sky130_fd_sc_hd__xnor2_2 _19521_ (.A(_17198_),
    .B(_17253_),
    .Y(_17264_));
 sky130_fd_sc_hd__xnor2_2 _19522_ (.A(_17188_),
    .B(_17264_),
    .Y(_17275_));
 sky130_fd_sc_hd__and3_2 _19523_ (.A(_17166_),
    .B(_17177_),
    .C(_17275_),
    .X(_17286_));
 sky130_fd_sc_hd__a21oi_2 _19524_ (.A1(_17166_),
    .A2(_17177_),
    .B1(_17275_),
    .Y(_17297_));
 sky130_fd_sc_hd__or2_2 _19525_ (.A(_17286_),
    .B(_17297_),
    .X(_17308_));
 sky130_fd_sc_hd__a21o_2 _19526_ (.A1(_16311_),
    .A2(_16432_),
    .B1(_17308_),
    .X(_17319_));
 sky130_fd_sc_hd__nand3_2 _19527_ (.A(_16311_),
    .B(_16432_),
    .C(_17308_),
    .Y(_17330_));
 sky130_fd_sc_hd__and2b_2 _19528_ (.A_N(_16640_),
    .B(_16629_),
    .X(_17341_));
 sky130_fd_sc_hd__or2b_2 _19529_ (.A(_16344_),
    .B_N(_16399_),
    .X(_17352_));
 sky130_fd_sc_hd__or2b_2 _19530_ (.A(_16333_),
    .B_N(_16410_),
    .X(_17363_));
 sky130_fd_sc_hd__and4_2 _19531_ (.A(iX[2]),
    .B(iX[3]),
    .C(iY[12]),
    .D(iY[13]),
    .X(_17374_));
 sky130_fd_sc_hd__a22oi_2 _19532_ (.A1(iX[3]),
    .A2(iY[12]),
    .B1(iY[13]),
    .B2(iX[2]),
    .Y(_17385_));
 sky130_fd_sc_hd__nor2_2 _19533_ (.A(_17374_),
    .B(_17385_),
    .Y(_17396_));
 sky130_fd_sc_hd__a21oi_2 _19534_ (.A1(iX[1]),
    .A2(iY[14]),
    .B1(_17396_),
    .Y(_17407_));
 sky130_fd_sc_hd__and3_2 _19535_ (.A(iX[1]),
    .B(iY[14]),
    .C(_17396_),
    .X(_17418_));
 sky130_fd_sc_hd__nor2_2 _19536_ (.A(_17407_),
    .B(_17418_),
    .Y(_17429_));
 sky130_fd_sc_hd__and4_2 _19537_ (.A(iX[5]),
    .B(iX[6]),
    .C(iY[9]),
    .D(iY[10]),
    .X(_17440_));
 sky130_fd_sc_hd__a22oi_2 _19538_ (.A1(iX[6]),
    .A2(iY[9]),
    .B1(iY[10]),
    .B2(iX[5]),
    .Y(_17451_));
 sky130_fd_sc_hd__nor2_2 _19539_ (.A(_17440_),
    .B(_17451_),
    .Y(_17462_));
 sky130_fd_sc_hd__nand2_2 _19540_ (.A(iX[4]),
    .B(iY[11]),
    .Y(_17473_));
 sky130_fd_sc_hd__xnor2_2 _19541_ (.A(_17462_),
    .B(_17473_),
    .Y(_17484_));
 sky130_fd_sc_hd__o21ba_2 _19542_ (.A1(_16596_),
    .A2(_16618_),
    .B1_N(_16585_),
    .X(_17495_));
 sky130_fd_sc_hd__xnor2_2 _19543_ (.A(_17484_),
    .B(_17495_),
    .Y(_17506_));
 sky130_fd_sc_hd__and2_2 _19544_ (.A(_17429_),
    .B(_17506_),
    .X(_17517_));
 sky130_fd_sc_hd__nor2_2 _19545_ (.A(_17429_),
    .B(_17506_),
    .Y(_17528_));
 sky130_fd_sc_hd__or2_2 _19546_ (.A(_17517_),
    .B(_17528_),
    .X(_17539_));
 sky130_fd_sc_hd__a21o_2 _19547_ (.A1(_17352_),
    .A2(_17363_),
    .B1(_17539_),
    .X(_17549_));
 sky130_fd_sc_hd__nand3_2 _19548_ (.A(_17352_),
    .B(_17363_),
    .C(_17539_),
    .Y(_17560_));
 sky130_fd_sc_hd__o211ai_2 _19549_ (.A1(_17341_),
    .A2(_16662_),
    .B1(_17549_),
    .C1(_17560_),
    .Y(_17571_));
 sky130_fd_sc_hd__a211o_2 _19550_ (.A1(_17549_),
    .A2(_17560_),
    .B1(_17341_),
    .C1(_16662_),
    .X(_17582_));
 sky130_fd_sc_hd__nand4_2 _19551_ (.A(_17319_),
    .B(_17330_),
    .C(_17571_),
    .D(_17582_),
    .Y(_17593_));
 sky130_fd_sc_hd__a22o_2 _19552_ (.A1(_17319_),
    .A2(_17330_),
    .B1(_17571_),
    .B2(_17582_),
    .X(_17604_));
 sky130_fd_sc_hd__o211ai_2 _19553_ (.A1(_16990_),
    .A2(_16750_),
    .B1(_17593_),
    .C1(_17604_),
    .Y(_17615_));
 sky130_fd_sc_hd__a211o_2 _19554_ (.A1(_17593_),
    .A2(_17604_),
    .B1(_16990_),
    .C1(_16750_),
    .X(_17626_));
 sky130_fd_sc_hd__o21ba_2 _19555_ (.A1(_16541_),
    .A2(_16563_),
    .B1_N(_16530_),
    .X(_17637_));
 sky130_fd_sc_hd__nand2_2 _19556_ (.A(iX[0]),
    .B(iY[15]),
    .Y(_17648_));
 sky130_fd_sc_hd__xnor2_2 _19557_ (.A(_17637_),
    .B(_17648_),
    .Y(_17659_));
 sky130_fd_sc_hd__a21o_2 _19558_ (.A1(_16695_),
    .A2(_16728_),
    .B1(_17659_),
    .X(_17670_));
 sky130_fd_sc_hd__nand3_2 _19559_ (.A(_16695_),
    .B(_16728_),
    .C(_17659_),
    .Y(_17681_));
 sky130_fd_sc_hd__and2_2 _19560_ (.A(_17670_),
    .B(_17681_),
    .X(_17692_));
 sky130_fd_sc_hd__a21oi_2 _19561_ (.A1(_17615_),
    .A2(_17626_),
    .B1(_17692_),
    .Y(_17703_));
 sky130_fd_sc_hd__and3_2 _19562_ (.A(_17615_),
    .B(_17626_),
    .C(_17692_),
    .X(_17714_));
 sky130_fd_sc_hd__nor2_2 _19563_ (.A(_17703_),
    .B(_17714_),
    .Y(_17725_));
 sky130_fd_sc_hd__a21bo_2 _19564_ (.A1(_16783_),
    .A2(_16826_),
    .B1_N(_16772_),
    .X(_17736_));
 sky130_fd_sc_hd__xnor2_2 _19565_ (.A(_17725_),
    .B(_17736_),
    .Y(_17747_));
 sky130_fd_sc_hd__xnor2_2 _19566_ (.A(_16805_),
    .B(_17747_),
    .Y(_17758_));
 sky130_fd_sc_hd__xor2_2 _19567_ (.A(_16979_),
    .B(_17758_),
    .X(_17769_));
 sky130_fd_sc_hd__inv_2 _19568_ (.A(_16892_),
    .Y(_17780_));
 sky130_fd_sc_hd__and2_2 _19569_ (.A(_16125_),
    .B(_17780_),
    .X(_17791_));
 sky130_fd_sc_hd__nor2_2 _19570_ (.A(_16914_),
    .B(_16903_),
    .Y(_17802_));
 sky130_fd_sc_hd__nor2_2 _19571_ (.A(_17791_),
    .B(_17802_),
    .Y(_17813_));
 sky130_fd_sc_hd__xnor2_2 _19572_ (.A(_17769_),
    .B(_17813_),
    .Y(_17824_));
 sky130_fd_sc_hd__xor2_2 _19573_ (.A(_16968_),
    .B(_17824_),
    .X(oO[15]));
 sky130_fd_sc_hd__a22oi_2 _19574_ (.A1(_17802_),
    .A2(_17769_),
    .B1(_17824_),
    .B2(_16968_),
    .Y(_17845_));
 sky130_fd_sc_hd__nor2_2 _19575_ (.A(_16979_),
    .B(_17758_),
    .Y(_17856_));
 sky130_fd_sc_hd__inv_2 _19576_ (.A(_17856_),
    .Y(_17867_));
 sky130_fd_sc_hd__a21boi_2 _19577_ (.A1(_17626_),
    .A2(_17692_),
    .B1_N(_17615_),
    .Y(_17878_));
 sky130_fd_sc_hd__or2b_2 _19578_ (.A(_17078_),
    .B_N(_17067_),
    .X(_17889_));
 sky130_fd_sc_hd__nand2_2 _19579_ (.A(_17089_),
    .B(_17144_),
    .Y(_17899_));
 sky130_fd_sc_hd__and4_2 _19580_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[15]),
    .D(iX[16]),
    .X(_17910_));
 sky130_fd_sc_hd__a22oi_2 _19581_ (.A1(iY[1]),
    .A2(iX[15]),
    .B1(iX[16]),
    .B2(iY[0]),
    .Y(_17921_));
 sky130_fd_sc_hd__nor2_2 _19582_ (.A(_17910_),
    .B(_17921_),
    .Y(_17932_));
 sky130_fd_sc_hd__nand2_2 _19583_ (.A(iY[2]),
    .B(iX[14]),
    .Y(_17943_));
 sky130_fd_sc_hd__xnor2_2 _19584_ (.A(_17932_),
    .B(_17943_),
    .Y(_17954_));
 sky130_fd_sc_hd__o21ba_2 _19585_ (.A1(_17034_),
    .A2(_17056_),
    .B1_N(_17023_),
    .X(_17965_));
 sky130_fd_sc_hd__xnor2_2 _19586_ (.A(_17954_),
    .B(_17965_),
    .Y(_17976_));
 sky130_fd_sc_hd__and4_2 _19587_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[12]),
    .D(iX[13]),
    .X(_17987_));
 sky130_fd_sc_hd__a22oi_2 _19588_ (.A1(iY[4]),
    .A2(iX[12]),
    .B1(iX[13]),
    .B2(iY[3]),
    .Y(_17998_));
 sky130_fd_sc_hd__nor2_2 _19589_ (.A(_17987_),
    .B(_17998_),
    .Y(_18009_));
 sky130_fd_sc_hd__nand2_2 _19590_ (.A(iY[5]),
    .B(iX[11]),
    .Y(_18020_));
 sky130_fd_sc_hd__xnor2_2 _19591_ (.A(_18009_),
    .B(_18020_),
    .Y(_18031_));
 sky130_fd_sc_hd__xnor2_2 _19592_ (.A(_17976_),
    .B(_18031_),
    .Y(_18042_));
 sky130_fd_sc_hd__a21o_2 _19593_ (.A1(_17889_),
    .A2(_17899_),
    .B1(_18042_),
    .X(_18053_));
 sky130_fd_sc_hd__nand3_2 _19594_ (.A(_17889_),
    .B(_17899_),
    .C(_18042_),
    .Y(_18064_));
 sky130_fd_sc_hd__o21ba_2 _19595_ (.A1(_17220_),
    .A2(_17242_),
    .B1_N(_17209_),
    .X(_18075_));
 sky130_fd_sc_hd__o21ba_2 _19596_ (.A1(_17111_),
    .A2(_17133_),
    .B1_N(_17100_),
    .X(_18086_));
 sky130_fd_sc_hd__and4_2 _19597_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[9]),
    .D(iX[10]),
    .X(_18097_));
 sky130_fd_sc_hd__a22oi_2 _19598_ (.A1(iY[7]),
    .A2(iX[9]),
    .B1(iX[10]),
    .B2(iY[6]),
    .Y(_18108_));
 sky130_fd_sc_hd__nor2_2 _19599_ (.A(_18097_),
    .B(_18108_),
    .Y(_18119_));
 sky130_fd_sc_hd__nand2_2 _19600_ (.A(iX[8]),
    .B(iY[8]),
    .Y(_18130_));
 sky130_fd_sc_hd__xnor2_2 _19601_ (.A(_18119_),
    .B(_18130_),
    .Y(_18141_));
 sky130_fd_sc_hd__xnor2_2 _19602_ (.A(_18086_),
    .B(_18141_),
    .Y(_18152_));
 sky130_fd_sc_hd__xnor2_2 _19603_ (.A(_18075_),
    .B(_18152_),
    .Y(_18163_));
 sky130_fd_sc_hd__nand3_2 _19604_ (.A(_18053_),
    .B(_18064_),
    .C(_18163_),
    .Y(_18174_));
 sky130_fd_sc_hd__a21o_2 _19605_ (.A1(_18053_),
    .A2(_18064_),
    .B1(_18163_),
    .X(_18185_));
 sky130_fd_sc_hd__a21bo_2 _19606_ (.A1(_17177_),
    .A2(_17275_),
    .B1_N(_17166_),
    .X(_18196_));
 sky130_fd_sc_hd__and3_2 _19607_ (.A(_18174_),
    .B(_18185_),
    .C(_18196_),
    .X(_18207_));
 sky130_fd_sc_hd__a21oi_2 _19608_ (.A1(_18174_),
    .A2(_18185_),
    .B1(_18196_),
    .Y(_18218_));
 sky130_fd_sc_hd__and2b_2 _19609_ (.A_N(_17495_),
    .B(_17484_),
    .X(_18229_));
 sky130_fd_sc_hd__or2b_2 _19610_ (.A(_17198_),
    .B_N(_17253_),
    .X(_18240_));
 sky130_fd_sc_hd__or2b_2 _19611_ (.A(_17188_),
    .B_N(_17264_),
    .X(_18251_));
 sky130_fd_sc_hd__and4_2 _19612_ (.A(iX[3]),
    .B(iX[4]),
    .C(iY[12]),
    .D(iY[13]),
    .X(_18262_));
 sky130_fd_sc_hd__a22o_2 _19613_ (.A1(iX[4]),
    .A2(iY[12]),
    .B1(iY[13]),
    .B2(iX[3]),
    .X(_18272_));
 sky130_fd_sc_hd__and2b_2 _19614_ (.A_N(_18262_),
    .B(_18272_),
    .X(_18283_));
 sky130_fd_sc_hd__nand2_2 _19615_ (.A(iX[2]),
    .B(iY[14]),
    .Y(_18294_));
 sky130_fd_sc_hd__xnor2_2 _19616_ (.A(_18283_),
    .B(_18294_),
    .Y(_18305_));
 sky130_fd_sc_hd__and4_2 _19617_ (.A(iX[6]),
    .B(iX[7]),
    .C(iY[9]),
    .D(iY[10]),
    .X(_18316_));
 sky130_fd_sc_hd__a22oi_2 _19618_ (.A1(iX[7]),
    .A2(iY[9]),
    .B1(iY[10]),
    .B2(iX[6]),
    .Y(_18327_));
 sky130_fd_sc_hd__nor2_2 _19619_ (.A(_18316_),
    .B(_18327_),
    .Y(_18338_));
 sky130_fd_sc_hd__nand2_2 _19620_ (.A(iX[5]),
    .B(iY[11]),
    .Y(_18349_));
 sky130_fd_sc_hd__xnor2_2 _19621_ (.A(_18338_),
    .B(_18349_),
    .Y(_18360_));
 sky130_fd_sc_hd__o21ba_2 _19622_ (.A1(_17451_),
    .A2(_17473_),
    .B1_N(_17440_),
    .X(_18371_));
 sky130_fd_sc_hd__xnor2_2 _19623_ (.A(_18360_),
    .B(_18371_),
    .Y(_18382_));
 sky130_fd_sc_hd__and2_2 _19624_ (.A(_18305_),
    .B(_18382_),
    .X(_18393_));
 sky130_fd_sc_hd__nor2_2 _19625_ (.A(_18305_),
    .B(_18382_),
    .Y(_18404_));
 sky130_fd_sc_hd__or2_2 _19626_ (.A(_18393_),
    .B(_18404_),
    .X(_18415_));
 sky130_fd_sc_hd__a21o_2 _19627_ (.A1(_18240_),
    .A2(_18251_),
    .B1(_18415_),
    .X(_18426_));
 sky130_fd_sc_hd__nand3_2 _19628_ (.A(_18240_),
    .B(_18251_),
    .C(_18415_),
    .Y(_18437_));
 sky130_fd_sc_hd__o211ai_2 _19629_ (.A1(_18229_),
    .A2(_17517_),
    .B1(_18426_),
    .C1(_18437_),
    .Y(_18448_));
 sky130_fd_sc_hd__a211o_2 _19630_ (.A1(_18426_),
    .A2(_18437_),
    .B1(_18229_),
    .C1(_17517_),
    .X(_18459_));
 sky130_fd_sc_hd__and4bb_2 _19631_ (.A_N(_18207_),
    .B_N(_18218_),
    .C(_18448_),
    .D(_18459_),
    .X(_18470_));
 sky130_fd_sc_hd__a2bb2oi_2 _19632_ (.A1_N(_18207_),
    .A2_N(_18218_),
    .B1(_18448_),
    .B2(_18459_),
    .Y(_18481_));
 sky130_fd_sc_hd__a211o_2 _19633_ (.A1(_17319_),
    .A2(_17593_),
    .B1(_18470_),
    .C1(_18481_),
    .X(_18492_));
 sky130_fd_sc_hd__o211ai_2 _19634_ (.A1(_18470_),
    .A2(_18481_),
    .B1(_17319_),
    .C1(_17593_),
    .Y(_18503_));
 sky130_fd_sc_hd__nand2_2 _19635_ (.A(_18492_),
    .B(_18503_),
    .Y(_18514_));
 sky130_fd_sc_hd__nor2_2 _19636_ (.A(_17637_),
    .B(_17648_),
    .Y(_18525_));
 sky130_fd_sc_hd__or2_2 _19637_ (.A(_17374_),
    .B(_17418_),
    .X(_18536_));
 sky130_fd_sc_hd__nand2_2 _19638_ (.A(iX[1]),
    .B(iY[16]),
    .Y(_18547_));
 sky130_fd_sc_hd__a22o_2 _19639_ (.A1(iX[1]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[0]),
    .X(_18558_));
 sky130_fd_sc_hd__o21ai_2 _19640_ (.A1(_17648_),
    .A2(_18547_),
    .B1(_18558_),
    .Y(_18569_));
 sky130_fd_sc_hd__xnor2_2 _19641_ (.A(_18536_),
    .B(_18569_),
    .Y(_18580_));
 sky130_fd_sc_hd__nand2_2 _19642_ (.A(_18525_),
    .B(_18580_),
    .Y(_18591_));
 sky130_fd_sc_hd__or2_2 _19643_ (.A(_18525_),
    .B(_18580_),
    .X(_18602_));
 sky130_fd_sc_hd__nand2_2 _19644_ (.A(_18591_),
    .B(_18602_),
    .Y(_18613_));
 sky130_fd_sc_hd__a21oi_2 _19645_ (.A1(_17549_),
    .A2(_17571_),
    .B1(_18613_),
    .Y(_18624_));
 sky130_fd_sc_hd__and3_2 _19646_ (.A(_17549_),
    .B(_17571_),
    .C(_18613_),
    .X(_18635_));
 sky130_fd_sc_hd__nor2_2 _19647_ (.A(_18624_),
    .B(_18635_),
    .Y(_18646_));
 sky130_fd_sc_hd__xnor2_2 _19648_ (.A(_18514_),
    .B(_18646_),
    .Y(_18657_));
 sky130_fd_sc_hd__or2b_2 _19649_ (.A(_17878_),
    .B_N(_18657_),
    .X(_18668_));
 sky130_fd_sc_hd__or2b_2 _19650_ (.A(_18657_),
    .B_N(_17878_),
    .X(_18678_));
 sky130_fd_sc_hd__nand2_2 _19651_ (.A(_18668_),
    .B(_18678_),
    .Y(_18689_));
 sky130_fd_sc_hd__xnor2_2 _19652_ (.A(_17670_),
    .B(_18689_),
    .Y(_18700_));
 sky130_fd_sc_hd__nand2_2 _19653_ (.A(_17725_),
    .B(_17736_),
    .Y(_18711_));
 sky130_fd_sc_hd__o21a_2 _19654_ (.A1(_16805_),
    .A2(_17747_),
    .B1(_18711_),
    .X(_18722_));
 sky130_fd_sc_hd__xnor2_2 _19655_ (.A(_18700_),
    .B(_18722_),
    .Y(_18733_));
 sky130_fd_sc_hd__and2_2 _19656_ (.A(_17791_),
    .B(_17769_),
    .X(_18744_));
 sky130_fd_sc_hd__xor2_2 _19657_ (.A(_18700_),
    .B(_18722_),
    .X(_18755_));
 sky130_fd_sc_hd__or3_2 _19658_ (.A(_17856_),
    .B(_18744_),
    .C(_18755_),
    .X(_18766_));
 sky130_fd_sc_hd__nand2_2 _19659_ (.A(_18744_),
    .B(_18755_),
    .Y(_18777_));
 sky130_fd_sc_hd__o211ai_2 _19660_ (.A1(_17867_),
    .A2(_18733_),
    .B1(_18766_),
    .C1(_18777_),
    .Y(_18788_));
 sky130_fd_sc_hd__xor2_2 _19661_ (.A(_17845_),
    .B(_18788_),
    .X(oO[16]));
 sky130_fd_sc_hd__nor2_2 _19662_ (.A(_17867_),
    .B(_18733_),
    .Y(_18809_));
 sky130_fd_sc_hd__or2_2 _19663_ (.A(_18700_),
    .B(_18722_),
    .X(_18820_));
 sky130_fd_sc_hd__or3_2 _19664_ (.A(_18514_),
    .B(_18624_),
    .C(_18635_),
    .X(_18831_));
 sky130_fd_sc_hd__or2b_2 _19665_ (.A(_17965_),
    .B_N(_17954_),
    .X(_18842_));
 sky130_fd_sc_hd__nand2_2 _19666_ (.A(_17976_),
    .B(_18031_),
    .Y(_18853_));
 sky130_fd_sc_hd__and4_2 _19667_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[16]),
    .D(iX[17]),
    .X(_18864_));
 sky130_fd_sc_hd__a22oi_2 _19668_ (.A1(iY[1]),
    .A2(iX[16]),
    .B1(iX[17]),
    .B2(iY[0]),
    .Y(_18875_));
 sky130_fd_sc_hd__nor2_2 _19669_ (.A(_18864_),
    .B(_18875_),
    .Y(_18886_));
 sky130_fd_sc_hd__nand2_2 _19670_ (.A(iY[2]),
    .B(iX[15]),
    .Y(_18897_));
 sky130_fd_sc_hd__xnor2_2 _19671_ (.A(_18886_),
    .B(_18897_),
    .Y(_18908_));
 sky130_fd_sc_hd__o21ba_2 _19672_ (.A1(_17921_),
    .A2(_17943_),
    .B1_N(_17910_),
    .X(_18919_));
 sky130_fd_sc_hd__xnor2_2 _19673_ (.A(_18908_),
    .B(_18919_),
    .Y(_00000_));
 sky130_fd_sc_hd__and4_2 _19674_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[13]),
    .D(iX[14]),
    .X(_00011_));
 sky130_fd_sc_hd__a22oi_2 _19675_ (.A1(iY[4]),
    .A2(iX[13]),
    .B1(iX[14]),
    .B2(iY[3]),
    .Y(_00022_));
 sky130_fd_sc_hd__nor2_2 _19676_ (.A(_00011_),
    .B(_00022_),
    .Y(_00033_));
 sky130_fd_sc_hd__nand2_2 _19677_ (.A(iY[5]),
    .B(iX[12]),
    .Y(_00044_));
 sky130_fd_sc_hd__xnor2_2 _19678_ (.A(_00033_),
    .B(_00044_),
    .Y(_00055_));
 sky130_fd_sc_hd__xnor2_2 _19679_ (.A(_00000_),
    .B(_00055_),
    .Y(_00066_));
 sky130_fd_sc_hd__a21o_2 _19680_ (.A1(_18842_),
    .A2(_18853_),
    .B1(_00066_),
    .X(_00077_));
 sky130_fd_sc_hd__nand3_2 _19681_ (.A(_18842_),
    .B(_18853_),
    .C(_00066_),
    .Y(_00088_));
 sky130_fd_sc_hd__o21ba_2 _19682_ (.A1(_18108_),
    .A2(_18130_),
    .B1_N(_18097_),
    .X(_00098_));
 sky130_fd_sc_hd__o21ba_2 _19683_ (.A1(_17998_),
    .A2(_18020_),
    .B1_N(_17987_),
    .X(_00109_));
 sky130_fd_sc_hd__and4_2 _19684_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[10]),
    .D(iX[11]),
    .X(_00120_));
 sky130_fd_sc_hd__a22oi_2 _19685_ (.A1(iY[7]),
    .A2(iX[10]),
    .B1(iX[11]),
    .B2(iY[6]),
    .Y(_00131_));
 sky130_fd_sc_hd__nor2_2 _19686_ (.A(_00120_),
    .B(_00131_),
    .Y(_00142_));
 sky130_fd_sc_hd__nand2_2 _19687_ (.A(iY[8]),
    .B(iX[9]),
    .Y(_00153_));
 sky130_fd_sc_hd__xnor2_2 _19688_ (.A(_00142_),
    .B(_00153_),
    .Y(_00164_));
 sky130_fd_sc_hd__xnor2_2 _19689_ (.A(_00109_),
    .B(_00164_),
    .Y(_00175_));
 sky130_fd_sc_hd__xnor2_2 _19690_ (.A(_00098_),
    .B(_00175_),
    .Y(_00186_));
 sky130_fd_sc_hd__nand3_2 _19691_ (.A(_00077_),
    .B(_00088_),
    .C(_00186_),
    .Y(_00197_));
 sky130_fd_sc_hd__a21o_2 _19692_ (.A1(_00077_),
    .A2(_00088_),
    .B1(_00186_),
    .X(_00208_));
 sky130_fd_sc_hd__nand2_2 _19693_ (.A(_18053_),
    .B(_18174_),
    .Y(_00219_));
 sky130_fd_sc_hd__and3_2 _19694_ (.A(_00197_),
    .B(_00208_),
    .C(_00219_),
    .X(_00230_));
 sky130_fd_sc_hd__a21oi_2 _19695_ (.A1(_00197_),
    .A2(_00208_),
    .B1(_00219_),
    .Y(_00241_));
 sky130_fd_sc_hd__and2b_2 _19696_ (.A_N(_18371_),
    .B(_18360_),
    .X(_00252_));
 sky130_fd_sc_hd__or2b_2 _19697_ (.A(_18086_),
    .B_N(_18141_),
    .X(_00263_));
 sky130_fd_sc_hd__or2b_2 _19698_ (.A(_18075_),
    .B_N(_18152_),
    .X(_00274_));
 sky130_fd_sc_hd__and4_2 _19699_ (.A(iX[4]),
    .B(iX[5]),
    .C(iY[12]),
    .D(iY[13]),
    .X(_00285_));
 sky130_fd_sc_hd__a22oi_2 _19700_ (.A1(iX[5]),
    .A2(iY[12]),
    .B1(iY[13]),
    .B2(iX[4]),
    .Y(_00296_));
 sky130_fd_sc_hd__nor2_2 _19701_ (.A(_00285_),
    .B(_00296_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand2_2 _19702_ (.A(iX[3]),
    .B(iY[14]),
    .Y(_00318_));
 sky130_fd_sc_hd__xnor2_2 _19703_ (.A(_00307_),
    .B(_00318_),
    .Y(_00329_));
 sky130_fd_sc_hd__and4_2 _19704_ (.A(iX[7]),
    .B(iX[8]),
    .C(iY[9]),
    .D(iY[10]),
    .X(_00340_));
 sky130_fd_sc_hd__a22oi_2 _19705_ (.A1(iX[8]),
    .A2(iY[9]),
    .B1(iY[10]),
    .B2(iX[7]),
    .Y(_00351_));
 sky130_fd_sc_hd__nor2_2 _19706_ (.A(_00340_),
    .B(_00351_),
    .Y(_00362_));
 sky130_fd_sc_hd__nand2_2 _19707_ (.A(iX[6]),
    .B(iY[11]),
    .Y(_00373_));
 sky130_fd_sc_hd__xnor2_2 _19708_ (.A(_00362_),
    .B(_00373_),
    .Y(_00384_));
 sky130_fd_sc_hd__o21ba_2 _19709_ (.A1(_18327_),
    .A2(_18349_),
    .B1_N(_18316_),
    .X(_00395_));
 sky130_fd_sc_hd__xnor2_2 _19710_ (.A(_00384_),
    .B(_00395_),
    .Y(_00406_));
 sky130_fd_sc_hd__and2_2 _19711_ (.A(_00329_),
    .B(_00406_),
    .X(_00417_));
 sky130_fd_sc_hd__nor2_2 _19712_ (.A(_00329_),
    .B(_00406_),
    .Y(_00428_));
 sky130_fd_sc_hd__or2_2 _19713_ (.A(_00417_),
    .B(_00428_),
    .X(_00439_));
 sky130_fd_sc_hd__a21o_2 _19714_ (.A1(_00263_),
    .A2(_00274_),
    .B1(_00439_),
    .X(_00450_));
 sky130_fd_sc_hd__nand3_2 _19715_ (.A(_00263_),
    .B(_00274_),
    .C(_00439_),
    .Y(_00461_));
 sky130_fd_sc_hd__o211ai_2 _19716_ (.A1(_00252_),
    .A2(_18393_),
    .B1(_00450_),
    .C1(_00461_),
    .Y(_00472_));
 sky130_fd_sc_hd__a211o_2 _19717_ (.A1(_00450_),
    .A2(_00461_),
    .B1(_00252_),
    .C1(_18393_),
    .X(_00483_));
 sky130_fd_sc_hd__and4bb_2 _19718_ (.A_N(_00230_),
    .B_N(_00241_),
    .C(_00472_),
    .D(_00483_),
    .X(_00493_));
 sky130_fd_sc_hd__a2bb2oi_2 _19719_ (.A1_N(_00230_),
    .A2_N(_00241_),
    .B1(_00472_),
    .B2(_00483_),
    .Y(_00504_));
 sky130_fd_sc_hd__nor2_2 _19720_ (.A(_00493_),
    .B(_00504_),
    .Y(_00515_));
 sky130_fd_sc_hd__nor2_2 _19721_ (.A(_18207_),
    .B(_18470_),
    .Y(_00526_));
 sky130_fd_sc_hd__xnor2_2 _19722_ (.A(_00515_),
    .B(_00526_),
    .Y(_00537_));
 sky130_fd_sc_hd__nand2_2 _19723_ (.A(_18426_),
    .B(_18448_),
    .Y(_00548_));
 sky130_fd_sc_hd__a31o_2 _19724_ (.A1(iX[2]),
    .A2(iY[14]),
    .A3(_18272_),
    .B1(_18262_),
    .X(_00559_));
 sky130_fd_sc_hd__nand2_2 _19725_ (.A(iX[2]),
    .B(iY[15]),
    .Y(_00570_));
 sky130_fd_sc_hd__and4_2 _19726_ (.A(iX[1]),
    .B(iX[2]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_00581_));
 sky130_fd_sc_hd__a21oi_2 _19727_ (.A1(_18547_),
    .A2(_00570_),
    .B1(_00581_),
    .Y(_00592_));
 sky130_fd_sc_hd__a21oi_2 _19728_ (.A1(iX[0]),
    .A2(iY[17]),
    .B1(_00592_),
    .Y(_00603_));
 sky130_fd_sc_hd__and3_2 _19729_ (.A(iX[0]),
    .B(iY[17]),
    .C(_00592_),
    .X(_00614_));
 sky130_fd_sc_hd__nor2_2 _19730_ (.A(_00603_),
    .B(_00614_),
    .Y(_00625_));
 sky130_fd_sc_hd__or2_2 _19731_ (.A(_00559_),
    .B(_00625_),
    .X(_00636_));
 sky130_fd_sc_hd__nand2_2 _19732_ (.A(_00559_),
    .B(_00625_),
    .Y(_00647_));
 sky130_fd_sc_hd__nand2_2 _19733_ (.A(_00636_),
    .B(_00647_),
    .Y(_00658_));
 sky130_fd_sc_hd__nor2_2 _19734_ (.A(_17648_),
    .B(_18547_),
    .Y(_00669_));
 sky130_fd_sc_hd__a21oi_2 _19735_ (.A1(_18536_),
    .A2(_18558_),
    .B1(_00669_),
    .Y(_00680_));
 sky130_fd_sc_hd__xor2_2 _19736_ (.A(_00658_),
    .B(_00680_),
    .X(_00691_));
 sky130_fd_sc_hd__xnor2_2 _19737_ (.A(_00548_),
    .B(_00691_),
    .Y(_00702_));
 sky130_fd_sc_hd__and2_2 _19738_ (.A(_18591_),
    .B(_00702_),
    .X(_00713_));
 sky130_fd_sc_hd__nor2_2 _19739_ (.A(_18591_),
    .B(_00702_),
    .Y(_00724_));
 sky130_fd_sc_hd__nor2_2 _19740_ (.A(_00713_),
    .B(_00724_),
    .Y(_00735_));
 sky130_fd_sc_hd__nor2_2 _19741_ (.A(_00537_),
    .B(_00735_),
    .Y(_00746_));
 sky130_fd_sc_hd__and2_2 _19742_ (.A(_00537_),
    .B(_00735_),
    .X(_00757_));
 sky130_fd_sc_hd__a211o_2 _19743_ (.A1(_18492_),
    .A2(_18831_),
    .B1(_00746_),
    .C1(_00757_),
    .X(_00768_));
 sky130_fd_sc_hd__o211ai_2 _19744_ (.A1(_00746_),
    .A2(_00757_),
    .B1(_18492_),
    .C1(_18831_),
    .Y(_00779_));
 sky130_fd_sc_hd__and3_2 _19745_ (.A(_18624_),
    .B(_00768_),
    .C(_00779_),
    .X(_00790_));
 sky130_fd_sc_hd__a21oi_2 _19746_ (.A1(_00768_),
    .A2(_00779_),
    .B1(_18624_),
    .Y(_00801_));
 sky130_fd_sc_hd__or2_2 _19747_ (.A(_00790_),
    .B(_00801_),
    .X(_00812_));
 sky130_fd_sc_hd__o21ai_2 _19748_ (.A1(_17670_),
    .A2(_18689_),
    .B1(_18668_),
    .Y(_00823_));
 sky130_fd_sc_hd__xor2_2 _19749_ (.A(_00812_),
    .B(_00823_),
    .X(_00834_));
 sky130_fd_sc_hd__xor2_2 _19750_ (.A(_18820_),
    .B(_00834_),
    .X(_00845_));
 sky130_fd_sc_hd__nor2_2 _19751_ (.A(_18809_),
    .B(_00845_),
    .Y(_00856_));
 sky130_fd_sc_hd__and2_2 _19752_ (.A(_18809_),
    .B(_00845_),
    .X(_00867_));
 sky130_fd_sc_hd__o221a_2 _19753_ (.A1(_17845_),
    .A2(_18788_),
    .B1(_00856_),
    .B2(_00867_),
    .C1(_18777_),
    .X(_00878_));
 sky130_fd_sc_hd__inv_2 _19754_ (.A(_00845_),
    .Y(_00889_));
 sky130_fd_sc_hd__o32a_2 _19755_ (.A1(_17845_),
    .A2(_18788_),
    .A3(_00889_),
    .B1(_00856_),
    .B2(_18777_),
    .X(_00899_));
 sky130_fd_sc_hd__and2b_2 _19756_ (.A_N(_00878_),
    .B(_00899_),
    .X(_00910_));
 sky130_fd_sc_hd__buf_1 _19757_ (.A(_00910_),
    .X(oO[17]));
 sky130_fd_sc_hd__nand2_2 _19758_ (.A(_18809_),
    .B(_00845_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand2_2 _19759_ (.A(_00931_),
    .B(_00899_),
    .Y(_00942_));
 sky130_fd_sc_hd__nor2_2 _19760_ (.A(_18820_),
    .B(_00834_),
    .Y(_00953_));
 sky130_fd_sc_hd__or3b_2 _19761_ (.A(_00790_),
    .B(_00801_),
    .C_N(_00823_),
    .X(_00964_));
 sky130_fd_sc_hd__and2b_2 _19762_ (.A_N(_00526_),
    .B(_00515_),
    .X(_00975_));
 sky130_fd_sc_hd__or2b_2 _19763_ (.A(_18919_),
    .B_N(_18908_),
    .X(_00986_));
 sky130_fd_sc_hd__nand2_2 _19764_ (.A(_00000_),
    .B(_00055_),
    .Y(_00997_));
 sky130_fd_sc_hd__and4_2 _19765_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[17]),
    .D(iX[18]),
    .X(_01008_));
 sky130_fd_sc_hd__a22oi_2 _19766_ (.A1(iY[1]),
    .A2(iX[17]),
    .B1(iX[18]),
    .B2(iY[0]),
    .Y(_01019_));
 sky130_fd_sc_hd__nor2_2 _19767_ (.A(_01008_),
    .B(_01019_),
    .Y(_01030_));
 sky130_fd_sc_hd__nand2_2 _19768_ (.A(iY[2]),
    .B(iX[16]),
    .Y(_01041_));
 sky130_fd_sc_hd__xnor2_2 _19769_ (.A(_01030_),
    .B(_01041_),
    .Y(_01052_));
 sky130_fd_sc_hd__o21ba_2 _19770_ (.A1(_18875_),
    .A2(_18897_),
    .B1_N(_18864_),
    .X(_01063_));
 sky130_fd_sc_hd__xnor2_2 _19771_ (.A(_01052_),
    .B(_01063_),
    .Y(_01074_));
 sky130_fd_sc_hd__and4_2 _19772_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[14]),
    .D(iX[15]),
    .X(_01085_));
 sky130_fd_sc_hd__a22oi_2 _19773_ (.A1(iY[4]),
    .A2(iX[14]),
    .B1(iX[15]),
    .B2(iY[3]),
    .Y(_01096_));
 sky130_fd_sc_hd__nor2_2 _19774_ (.A(_01085_),
    .B(_01096_),
    .Y(_01107_));
 sky130_fd_sc_hd__nand2_2 _19775_ (.A(iY[5]),
    .B(iX[13]),
    .Y(_01118_));
 sky130_fd_sc_hd__xnor2_2 _19776_ (.A(_01107_),
    .B(_01118_),
    .Y(_01129_));
 sky130_fd_sc_hd__xnor2_2 _19777_ (.A(_01074_),
    .B(_01129_),
    .Y(_01140_));
 sky130_fd_sc_hd__a21o_2 _19778_ (.A1(_00986_),
    .A2(_00997_),
    .B1(_01140_),
    .X(_01151_));
 sky130_fd_sc_hd__nand3_2 _19779_ (.A(_00986_),
    .B(_00997_),
    .C(_01140_),
    .Y(_01162_));
 sky130_fd_sc_hd__o21ba_2 _19780_ (.A1(_00131_),
    .A2(_00153_),
    .B1_N(_00120_),
    .X(_01173_));
 sky130_fd_sc_hd__o21ba_2 _19781_ (.A1(_00022_),
    .A2(_00044_),
    .B1_N(_00011_),
    .X(_01184_));
 sky130_fd_sc_hd__and4_2 _19782_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[11]),
    .D(iX[12]),
    .X(_01195_));
 sky130_fd_sc_hd__a22oi_2 _19783_ (.A1(iY[7]),
    .A2(iX[11]),
    .B1(iX[12]),
    .B2(iY[6]),
    .Y(_01206_));
 sky130_fd_sc_hd__nor2_2 _19784_ (.A(_01195_),
    .B(_01206_),
    .Y(_01217_));
 sky130_fd_sc_hd__nand2_2 _19785_ (.A(iY[8]),
    .B(iX[10]),
    .Y(_01228_));
 sky130_fd_sc_hd__xnor2_2 _19786_ (.A(_01217_),
    .B(_01228_),
    .Y(_01239_));
 sky130_fd_sc_hd__xnor2_2 _19787_ (.A(_01184_),
    .B(_01239_),
    .Y(_01250_));
 sky130_fd_sc_hd__xnor2_2 _19788_ (.A(_01173_),
    .B(_01250_),
    .Y(_01261_));
 sky130_fd_sc_hd__nand3_2 _19789_ (.A(_01151_),
    .B(_01162_),
    .C(_01261_),
    .Y(_01272_));
 sky130_fd_sc_hd__a21o_2 _19790_ (.A1(_01151_),
    .A2(_01162_),
    .B1(_01261_),
    .X(_01283_));
 sky130_fd_sc_hd__nand2_2 _19791_ (.A(_01272_),
    .B(_01283_),
    .Y(_01294_));
 sky130_fd_sc_hd__nand2_2 _19792_ (.A(_00077_),
    .B(_00197_),
    .Y(_01305_));
 sky130_fd_sc_hd__xnor2_2 _19793_ (.A(_01294_),
    .B(_01305_),
    .Y(_01316_));
 sky130_fd_sc_hd__and2b_2 _19794_ (.A_N(_00395_),
    .B(_00384_),
    .X(_01326_));
 sky130_fd_sc_hd__or2b_2 _19795_ (.A(_00109_),
    .B_N(_00164_),
    .X(_01337_));
 sky130_fd_sc_hd__or2b_2 _19796_ (.A(_00098_),
    .B_N(_00175_),
    .X(_01348_));
 sky130_fd_sc_hd__and4_2 _19797_ (.A(iX[5]),
    .B(iX[6]),
    .C(iY[12]),
    .D(iY[13]),
    .X(_01359_));
 sky130_fd_sc_hd__a22oi_2 _19798_ (.A1(iX[6]),
    .A2(iY[12]),
    .B1(iY[13]),
    .B2(iX[5]),
    .Y(_01370_));
 sky130_fd_sc_hd__nor2_2 _19799_ (.A(_01359_),
    .B(_01370_),
    .Y(_01381_));
 sky130_fd_sc_hd__nand2_2 _19800_ (.A(iX[4]),
    .B(iY[14]),
    .Y(_01392_));
 sky130_fd_sc_hd__xnor2_2 _19801_ (.A(_01381_),
    .B(_01392_),
    .Y(_01403_));
 sky130_fd_sc_hd__and4_2 _19802_ (.A(iX[8]),
    .B(iX[9]),
    .C(iY[9]),
    .D(iY[10]),
    .X(_01414_));
 sky130_fd_sc_hd__a22oi_2 _19803_ (.A1(iX[9]),
    .A2(iY[9]),
    .B1(iY[10]),
    .B2(iX[8]),
    .Y(_01425_));
 sky130_fd_sc_hd__nor2_2 _19804_ (.A(_01414_),
    .B(_01425_),
    .Y(_01436_));
 sky130_fd_sc_hd__nand2_2 _19805_ (.A(iX[7]),
    .B(iY[11]),
    .Y(_01447_));
 sky130_fd_sc_hd__xnor2_2 _19806_ (.A(_01436_),
    .B(_01447_),
    .Y(_01458_));
 sky130_fd_sc_hd__o21ba_2 _19807_ (.A1(_00351_),
    .A2(_00373_),
    .B1_N(_00340_),
    .X(_01469_));
 sky130_fd_sc_hd__xnor2_2 _19808_ (.A(_01458_),
    .B(_01469_),
    .Y(_01480_));
 sky130_fd_sc_hd__and2_2 _19809_ (.A(_01403_),
    .B(_01480_),
    .X(_01491_));
 sky130_fd_sc_hd__nor2_2 _19810_ (.A(_01403_),
    .B(_01480_),
    .Y(_01502_));
 sky130_fd_sc_hd__or2_2 _19811_ (.A(_01491_),
    .B(_01502_),
    .X(_01513_));
 sky130_fd_sc_hd__a21o_2 _19812_ (.A1(_01337_),
    .A2(_01348_),
    .B1(_01513_),
    .X(_01524_));
 sky130_fd_sc_hd__nand3_2 _19813_ (.A(_01337_),
    .B(_01348_),
    .C(_01513_),
    .Y(_01535_));
 sky130_fd_sc_hd__o211ai_2 _19814_ (.A1(_01326_),
    .A2(_00417_),
    .B1(_01524_),
    .C1(_01535_),
    .Y(_01546_));
 sky130_fd_sc_hd__a211o_2 _19815_ (.A1(_01524_),
    .A2(_01535_),
    .B1(_01326_),
    .C1(_00417_),
    .X(_01557_));
 sky130_fd_sc_hd__and3_2 _19816_ (.A(_01316_),
    .B(_01546_),
    .C(_01557_),
    .X(_01568_));
 sky130_fd_sc_hd__inv_2 _19817_ (.A(_01568_),
    .Y(_01579_));
 sky130_fd_sc_hd__a21o_2 _19818_ (.A1(_01546_),
    .A2(_01557_),
    .B1(_01316_),
    .X(_01590_));
 sky130_fd_sc_hd__o211a_2 _19819_ (.A1(_00230_),
    .A2(_00493_),
    .B1(_01579_),
    .C1(_01590_),
    .X(_01601_));
 sky130_fd_sc_hd__a211oi_2 _19820_ (.A1(_01579_),
    .A2(_01590_),
    .B1(_00230_),
    .C1(_00493_),
    .Y(_01612_));
 sky130_fd_sc_hd__and4b_2 _19821_ (.A_N(_18569_),
    .B(_00636_),
    .C(_00647_),
    .D(_18536_),
    .X(_01623_));
 sky130_fd_sc_hd__nand2_2 _19822_ (.A(_00450_),
    .B(_00472_),
    .Y(_01634_));
 sky130_fd_sc_hd__o21ba_2 _19823_ (.A1(_00296_),
    .A2(_00318_),
    .B1_N(_00285_),
    .X(_01645_));
 sky130_fd_sc_hd__nand4_2 _19824_ (.A(iX[2]),
    .B(iX[3]),
    .C(iY[15]),
    .D(iY[16]),
    .Y(_01656_));
 sky130_fd_sc_hd__a22o_2 _19825_ (.A1(iX[3]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[2]),
    .X(_01667_));
 sky130_fd_sc_hd__and2_2 _19826_ (.A(iX[1]),
    .B(iY[17]),
    .X(_01678_));
 sky130_fd_sc_hd__a21oi_2 _19827_ (.A1(_01656_),
    .A2(_01667_),
    .B1(_01678_),
    .Y(_01689_));
 sky130_fd_sc_hd__and3_2 _19828_ (.A(_01656_),
    .B(_01667_),
    .C(_01678_),
    .X(_01700_));
 sky130_fd_sc_hd__nor2_2 _19829_ (.A(_01689_),
    .B(_01700_),
    .Y(_01711_));
 sky130_fd_sc_hd__xnor2_2 _19830_ (.A(_01645_),
    .B(_01711_),
    .Y(_01721_));
 sky130_fd_sc_hd__or3_2 _19831_ (.A(_00581_),
    .B(_00614_),
    .C(_01721_),
    .X(_01732_));
 sky130_fd_sc_hd__o21ai_2 _19832_ (.A1(_00581_),
    .A2(_00614_),
    .B1(_01721_),
    .Y(_01743_));
 sky130_fd_sc_hd__nand2_2 _19833_ (.A(_01732_),
    .B(_01743_),
    .Y(_01754_));
 sky130_fd_sc_hd__a21boi_2 _19834_ (.A1(_00669_),
    .A2(_00636_),
    .B1_N(_00647_),
    .Y(_01765_));
 sky130_fd_sc_hd__and2_2 _19835_ (.A(_01754_),
    .B(_01765_),
    .X(_01776_));
 sky130_fd_sc_hd__nor2_2 _19836_ (.A(_01754_),
    .B(_01765_),
    .Y(_01787_));
 sky130_fd_sc_hd__nor2_2 _19837_ (.A(_01776_),
    .B(_01787_),
    .Y(_01798_));
 sky130_fd_sc_hd__and2_2 _19838_ (.A(iX[0]),
    .B(iY[18]),
    .X(_01809_));
 sky130_fd_sc_hd__nor2_2 _19839_ (.A(_01798_),
    .B(_01809_),
    .Y(_01820_));
 sky130_fd_sc_hd__and2_2 _19840_ (.A(_01798_),
    .B(_01809_),
    .X(_01831_));
 sky130_fd_sc_hd__or2_2 _19841_ (.A(_01820_),
    .B(_01831_),
    .X(_01842_));
 sky130_fd_sc_hd__xor2_2 _19842_ (.A(_01634_),
    .B(_01842_),
    .X(_01853_));
 sky130_fd_sc_hd__xor2_2 _19843_ (.A(_01623_),
    .B(_01853_),
    .X(_01864_));
 sky130_fd_sc_hd__o21ai_2 _19844_ (.A1(_01601_),
    .A2(_01612_),
    .B1(_01864_),
    .Y(_01875_));
 sky130_fd_sc_hd__or3_2 _19845_ (.A(_01601_),
    .B(_01612_),
    .C(_01864_),
    .X(_01886_));
 sky130_fd_sc_hd__o211a_2 _19846_ (.A1(_00975_),
    .A2(_00757_),
    .B1(_01875_),
    .C1(_01886_),
    .X(_01897_));
 sky130_fd_sc_hd__a211oi_2 _19847_ (.A1(_01875_),
    .A2(_01886_),
    .B1(_00975_),
    .C1(_00757_),
    .Y(_01908_));
 sky130_fd_sc_hd__or2_2 _19848_ (.A(_01897_),
    .B(_01908_),
    .X(_01919_));
 sky130_fd_sc_hd__a21oi_2 _19849_ (.A1(_00548_),
    .A2(_00691_),
    .B1(_00724_),
    .Y(_01930_));
 sky130_fd_sc_hd__xnor2_2 _19850_ (.A(_01919_),
    .B(_01930_),
    .Y(_01941_));
 sky130_fd_sc_hd__a21bo_2 _19851_ (.A1(_18624_),
    .A2(_00779_),
    .B1_N(_00768_),
    .X(_01952_));
 sky130_fd_sc_hd__xnor2_2 _19852_ (.A(_01941_),
    .B(_01952_),
    .Y(_01963_));
 sky130_fd_sc_hd__xor2_2 _19853_ (.A(_00964_),
    .B(_01963_),
    .X(_01974_));
 sky130_fd_sc_hd__xnor2_2 _19854_ (.A(_00953_),
    .B(_01974_),
    .Y(_01985_));
 sky130_fd_sc_hd__xor2_2 _19855_ (.A(_00942_),
    .B(_01985_),
    .X(oO[18]));
 sky130_fd_sc_hd__or2b_2 _19856_ (.A(_00964_),
    .B_N(_01963_),
    .X(_02006_));
 sky130_fd_sc_hd__and2b_2 _19857_ (.A_N(_01941_),
    .B(_01952_),
    .X(_02017_));
 sky130_fd_sc_hd__nor3_2 _19858_ (.A(_01601_),
    .B(_01612_),
    .C(_01864_),
    .Y(_02028_));
 sky130_fd_sc_hd__and2b_2 _19859_ (.A_N(_01469_),
    .B(_01458_),
    .X(_02039_));
 sky130_fd_sc_hd__or2b_2 _19860_ (.A(_01184_),
    .B_N(_01239_),
    .X(_02050_));
 sky130_fd_sc_hd__or2b_2 _19861_ (.A(_01173_),
    .B_N(_01250_),
    .X(_02061_));
 sky130_fd_sc_hd__and4_2 _19862_ (.A(iX[6]),
    .B(iX[7]),
    .C(iY[12]),
    .D(iY[13]),
    .X(_02072_));
 sky130_fd_sc_hd__a22oi_2 _19863_ (.A1(iX[7]),
    .A2(iY[12]),
    .B1(iY[13]),
    .B2(iX[6]),
    .Y(_02083_));
 sky130_fd_sc_hd__nor2_2 _19864_ (.A(_02072_),
    .B(_02083_),
    .Y(_02094_));
 sky130_fd_sc_hd__nand2_2 _19865_ (.A(iX[5]),
    .B(iY[14]),
    .Y(_02105_));
 sky130_fd_sc_hd__xnor2_2 _19866_ (.A(_02094_),
    .B(_02105_),
    .Y(_02115_));
 sky130_fd_sc_hd__and4_2 _19867_ (.A(iX[9]),
    .B(iY[9]),
    .C(iX[10]),
    .D(iY[10]),
    .X(_02126_));
 sky130_fd_sc_hd__a22oi_2 _19868_ (.A1(iY[9]),
    .A2(iX[10]),
    .B1(iY[10]),
    .B2(iX[9]),
    .Y(_02137_));
 sky130_fd_sc_hd__nor2_2 _19869_ (.A(_02126_),
    .B(_02137_),
    .Y(_02148_));
 sky130_fd_sc_hd__nand2_2 _19870_ (.A(iX[8]),
    .B(iY[11]),
    .Y(_02159_));
 sky130_fd_sc_hd__xnor2_2 _19871_ (.A(_02148_),
    .B(_02159_),
    .Y(_02170_));
 sky130_fd_sc_hd__o21ba_2 _19872_ (.A1(_01425_),
    .A2(_01447_),
    .B1_N(_01414_),
    .X(_02181_));
 sky130_fd_sc_hd__xnor2_2 _19873_ (.A(_02170_),
    .B(_02181_),
    .Y(_02192_));
 sky130_fd_sc_hd__and2_2 _19874_ (.A(_02115_),
    .B(_02192_),
    .X(_02203_));
 sky130_fd_sc_hd__nor2_2 _19875_ (.A(_02115_),
    .B(_02192_),
    .Y(_02214_));
 sky130_fd_sc_hd__or2_2 _19876_ (.A(_02203_),
    .B(_02214_),
    .X(_02225_));
 sky130_fd_sc_hd__a21o_2 _19877_ (.A1(_02050_),
    .A2(_02061_),
    .B1(_02225_),
    .X(_02236_));
 sky130_fd_sc_hd__nand3_2 _19878_ (.A(_02050_),
    .B(_02061_),
    .C(_02225_),
    .Y(_02247_));
 sky130_fd_sc_hd__o211ai_2 _19879_ (.A1(_02039_),
    .A2(_01491_),
    .B1(_02236_),
    .C1(_02247_),
    .Y(_02258_));
 sky130_fd_sc_hd__a211o_2 _19880_ (.A1(_02236_),
    .A2(_02247_),
    .B1(_02039_),
    .C1(_01491_),
    .X(_02269_));
 sky130_fd_sc_hd__or2b_2 _19881_ (.A(_01063_),
    .B_N(_01052_),
    .X(_02280_));
 sky130_fd_sc_hd__nand2_2 _19882_ (.A(_01074_),
    .B(_01129_),
    .Y(_02291_));
 sky130_fd_sc_hd__and4_2 _19883_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[18]),
    .D(iX[19]),
    .X(_02302_));
 sky130_fd_sc_hd__a22oi_2 _19884_ (.A1(iY[1]),
    .A2(iX[18]),
    .B1(iX[19]),
    .B2(iY[0]),
    .Y(_02313_));
 sky130_fd_sc_hd__nor2_2 _19885_ (.A(_02302_),
    .B(_02313_),
    .Y(_02324_));
 sky130_fd_sc_hd__nand2_2 _19886_ (.A(iY[2]),
    .B(iX[17]),
    .Y(_02335_));
 sky130_fd_sc_hd__xnor2_2 _19887_ (.A(_02324_),
    .B(_02335_),
    .Y(_02346_));
 sky130_fd_sc_hd__o21ba_2 _19888_ (.A1(_01019_),
    .A2(_01041_),
    .B1_N(_01008_),
    .X(_02357_));
 sky130_fd_sc_hd__xnor2_2 _19889_ (.A(_02346_),
    .B(_02357_),
    .Y(_02368_));
 sky130_fd_sc_hd__and4_2 _19890_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[15]),
    .D(iX[16]),
    .X(_02379_));
 sky130_fd_sc_hd__a22oi_2 _19891_ (.A1(iY[4]),
    .A2(iX[15]),
    .B1(iX[16]),
    .B2(iY[3]),
    .Y(_02390_));
 sky130_fd_sc_hd__nor2_2 _19892_ (.A(_02379_),
    .B(_02390_),
    .Y(_02401_));
 sky130_fd_sc_hd__nand2_2 _19893_ (.A(iY[5]),
    .B(iX[14]),
    .Y(_02412_));
 sky130_fd_sc_hd__xnor2_2 _19894_ (.A(_02401_),
    .B(_02412_),
    .Y(_02423_));
 sky130_fd_sc_hd__xnor2_2 _19895_ (.A(_02368_),
    .B(_02423_),
    .Y(_02434_));
 sky130_fd_sc_hd__a21o_2 _19896_ (.A1(_02280_),
    .A2(_02291_),
    .B1(_02434_),
    .X(_02445_));
 sky130_fd_sc_hd__nand3_2 _19897_ (.A(_02280_),
    .B(_02291_),
    .C(_02434_),
    .Y(_02456_));
 sky130_fd_sc_hd__o21ba_2 _19898_ (.A1(_01206_),
    .A2(_01228_),
    .B1_N(_01195_),
    .X(_02467_));
 sky130_fd_sc_hd__o21ba_2 _19899_ (.A1(_01096_),
    .A2(_01118_),
    .B1_N(_01085_),
    .X(_02478_));
 sky130_fd_sc_hd__and4_2 _19900_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[12]),
    .D(iX[13]),
    .X(_02489_));
 sky130_fd_sc_hd__a22oi_2 _19901_ (.A1(iY[7]),
    .A2(iX[12]),
    .B1(iX[13]),
    .B2(iY[6]),
    .Y(_02500_));
 sky130_fd_sc_hd__nor2_2 _19902_ (.A(_02489_),
    .B(_02500_),
    .Y(_02511_));
 sky130_fd_sc_hd__nand2_2 _19903_ (.A(iY[8]),
    .B(iX[11]),
    .Y(_02521_));
 sky130_fd_sc_hd__xnor2_2 _19904_ (.A(_02511_),
    .B(_02521_),
    .Y(_02532_));
 sky130_fd_sc_hd__xnor2_2 _19905_ (.A(_02478_),
    .B(_02532_),
    .Y(_02543_));
 sky130_fd_sc_hd__xnor2_2 _19906_ (.A(_02467_),
    .B(_02543_),
    .Y(_02554_));
 sky130_fd_sc_hd__nand3_2 _19907_ (.A(_02445_),
    .B(_02456_),
    .C(_02554_),
    .Y(_02565_));
 sky130_fd_sc_hd__a21o_2 _19908_ (.A1(_02445_),
    .A2(_02456_),
    .B1(_02554_),
    .X(_02576_));
 sky130_fd_sc_hd__nand2_2 _19909_ (.A(_02565_),
    .B(_02576_),
    .Y(_02587_));
 sky130_fd_sc_hd__nand2_2 _19910_ (.A(_01151_),
    .B(_01272_),
    .Y(_02598_));
 sky130_fd_sc_hd__xnor2_2 _19911_ (.A(_02587_),
    .B(_02598_),
    .Y(_02609_));
 sky130_fd_sc_hd__a21oi_2 _19912_ (.A1(_02258_),
    .A2(_02269_),
    .B1(_02609_),
    .Y(_02620_));
 sky130_fd_sc_hd__and3_2 _19913_ (.A(_02609_),
    .B(_02258_),
    .C(_02269_),
    .X(_02631_));
 sky130_fd_sc_hd__a31oi_2 _19914_ (.A1(_01272_),
    .A2(_01283_),
    .A3(_01305_),
    .B1(_01568_),
    .Y(_02642_));
 sky130_fd_sc_hd__or3_2 _19915_ (.A(_02620_),
    .B(_02631_),
    .C(_02642_),
    .X(_02653_));
 sky130_fd_sc_hd__o21ai_2 _19916_ (.A1(_02620_),
    .A2(_02631_),
    .B1(_02642_),
    .Y(_02664_));
 sky130_fd_sc_hd__nand2_2 _19917_ (.A(_01524_),
    .B(_01546_),
    .Y(_02675_));
 sky130_fd_sc_hd__a22oi_2 _19918_ (.A1(iX[1]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[0]),
    .Y(_02686_));
 sky130_fd_sc_hd__and3_2 _19919_ (.A(iX[1]),
    .B(iY[19]),
    .C(_01809_),
    .X(_02697_));
 sky130_fd_sc_hd__or3_2 _19920_ (.A(_01645_),
    .B(_01689_),
    .C(_01700_),
    .X(_02708_));
 sky130_fd_sc_hd__and4_2 _19921_ (.A(iX[2]),
    .B(iX[3]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_02719_));
 sky130_fd_sc_hd__o21ba_2 _19922_ (.A1(_01370_),
    .A2(_01392_),
    .B1_N(_01359_),
    .X(_02730_));
 sky130_fd_sc_hd__and4_2 _19923_ (.A(iX[3]),
    .B(iX[4]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_02741_));
 sky130_fd_sc_hd__a22oi_2 _19924_ (.A1(iX[4]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[3]),
    .Y(_02752_));
 sky130_fd_sc_hd__nor2_2 _19925_ (.A(_02741_),
    .B(_02752_),
    .Y(_02763_));
 sky130_fd_sc_hd__nand2_2 _19926_ (.A(iX[2]),
    .B(iY[17]),
    .Y(_02774_));
 sky130_fd_sc_hd__xnor2_2 _19927_ (.A(_02763_),
    .B(_02774_),
    .Y(_02785_));
 sky130_fd_sc_hd__xnor2_2 _19928_ (.A(_02730_),
    .B(_02785_),
    .Y(_02796_));
 sky130_fd_sc_hd__o21ai_2 _19929_ (.A1(_02719_),
    .A2(_01700_),
    .B1(_02796_),
    .Y(_02807_));
 sky130_fd_sc_hd__or3_2 _19930_ (.A(_02719_),
    .B(_01700_),
    .C(_02796_),
    .X(_02818_));
 sky130_fd_sc_hd__nand2_2 _19931_ (.A(_02807_),
    .B(_02818_),
    .Y(_02829_));
 sky130_fd_sc_hd__a21o_2 _19932_ (.A1(_02708_),
    .A2(_01743_),
    .B1(_02829_),
    .X(_02840_));
 sky130_fd_sc_hd__nand3_2 _19933_ (.A(_02708_),
    .B(_01743_),
    .C(_02829_),
    .Y(_02851_));
 sky130_fd_sc_hd__nand2_2 _19934_ (.A(_02840_),
    .B(_02851_),
    .Y(_02862_));
 sky130_fd_sc_hd__or3_2 _19935_ (.A(_02686_),
    .B(_02697_),
    .C(_02862_),
    .X(_02873_));
 sky130_fd_sc_hd__o21ai_2 _19936_ (.A1(_02686_),
    .A2(_02697_),
    .B1(_02862_),
    .Y(_02884_));
 sky130_fd_sc_hd__and3_2 _19937_ (.A(_02675_),
    .B(_02873_),
    .C(_02884_),
    .X(_02895_));
 sky130_fd_sc_hd__a21oi_2 _19938_ (.A1(_02873_),
    .A2(_02884_),
    .B1(_02675_),
    .Y(_02906_));
 sky130_fd_sc_hd__nor2_2 _19939_ (.A(_02895_),
    .B(_02906_),
    .Y(_02916_));
 sky130_fd_sc_hd__o21ai_2 _19940_ (.A1(_01787_),
    .A2(_01831_),
    .B1(_02916_),
    .Y(_02927_));
 sky130_fd_sc_hd__or3_2 _19941_ (.A(_01787_),
    .B(_01831_),
    .C(_02916_),
    .X(_02938_));
 sky130_fd_sc_hd__nand4_2 _19942_ (.A(_02653_),
    .B(_02664_),
    .C(_02927_),
    .D(_02938_),
    .Y(_02949_));
 sky130_fd_sc_hd__a22o_2 _19943_ (.A1(_02653_),
    .A2(_02664_),
    .B1(_02927_),
    .B2(_02938_),
    .X(_02960_));
 sky130_fd_sc_hd__o211a_2 _19944_ (.A1(_01601_),
    .A2(_02028_),
    .B1(_02949_),
    .C1(_02960_),
    .X(_02971_));
 sky130_fd_sc_hd__a211o_2 _19945_ (.A1(_02949_),
    .A2(_02960_),
    .B1(_01601_),
    .C1(_02028_),
    .X(_02982_));
 sky130_fd_sc_hd__and2b_2 _19946_ (.A_N(_02971_),
    .B(_02982_),
    .X(_02993_));
 sky130_fd_sc_hd__inv_2 _19947_ (.A(_01853_),
    .Y(_03004_));
 sky130_fd_sc_hd__and2b_2 _19948_ (.A_N(_01842_),
    .B(_01634_),
    .X(_03015_));
 sky130_fd_sc_hd__a21o_2 _19949_ (.A1(_01623_),
    .A2(_03004_),
    .B1(_03015_),
    .X(_03026_));
 sky130_fd_sc_hd__xnor2_2 _19950_ (.A(_02993_),
    .B(_03026_),
    .Y(_03037_));
 sky130_fd_sc_hd__o21ba_2 _19951_ (.A1(_01919_),
    .A2(_01930_),
    .B1_N(_01897_),
    .X(_03048_));
 sky130_fd_sc_hd__xor2_2 _19952_ (.A(_03037_),
    .B(_03048_),
    .X(_03059_));
 sky130_fd_sc_hd__xnor2_2 _19953_ (.A(_02017_),
    .B(_03059_),
    .Y(_03070_));
 sky130_fd_sc_hd__xor2_2 _19954_ (.A(_02006_),
    .B(_03070_),
    .X(_03081_));
 sky130_fd_sc_hd__or3_2 _19955_ (.A(_18820_),
    .B(_00834_),
    .C(_01974_),
    .X(_03092_));
 sky130_fd_sc_hd__a21bo_2 _19956_ (.A1(_00942_),
    .A2(_01985_),
    .B1_N(_03092_),
    .X(_03103_));
 sky130_fd_sc_hd__xnor2_2 _19957_ (.A(_03081_),
    .B(_03103_),
    .Y(_03114_));
 sky130_fd_sc_hd__inv_2 _19958_ (.A(_03114_),
    .Y(oO[19]));
 sky130_fd_sc_hd__nand2_2 _19959_ (.A(_01985_),
    .B(_03081_),
    .Y(_03135_));
 sky130_fd_sc_hd__a21o_2 _19960_ (.A1(_00931_),
    .A2(_00899_),
    .B1(_03135_),
    .X(_03146_));
 sky130_fd_sc_hd__a21o_2 _19961_ (.A1(_02006_),
    .A2(_03092_),
    .B1(_03070_),
    .X(_03157_));
 sky130_fd_sc_hd__nand2_2 _19962_ (.A(_03146_),
    .B(_03157_),
    .Y(_03168_));
 sky130_fd_sc_hd__and3_2 _19963_ (.A(_02565_),
    .B(_02576_),
    .C(_02598_),
    .X(_03179_));
 sky130_fd_sc_hd__or2b_2 _19964_ (.A(_02357_),
    .B_N(_02346_),
    .X(_03190_));
 sky130_fd_sc_hd__nand2_2 _19965_ (.A(_02368_),
    .B(_02423_),
    .Y(_03201_));
 sky130_fd_sc_hd__and4_2 _19966_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[19]),
    .D(iX[20]),
    .X(_03212_));
 sky130_fd_sc_hd__a22oi_2 _19967_ (.A1(iY[1]),
    .A2(iX[19]),
    .B1(iX[20]),
    .B2(iY[0]),
    .Y(_03223_));
 sky130_fd_sc_hd__nor2_2 _19968_ (.A(_03212_),
    .B(_03223_),
    .Y(_03234_));
 sky130_fd_sc_hd__nand2_2 _19969_ (.A(iY[2]),
    .B(iX[18]),
    .Y(_03245_));
 sky130_fd_sc_hd__xnor2_2 _19970_ (.A(_03234_),
    .B(_03245_),
    .Y(_03256_));
 sky130_fd_sc_hd__o21ba_2 _19971_ (.A1(_02313_),
    .A2(_02335_),
    .B1_N(_02302_),
    .X(_03267_));
 sky130_fd_sc_hd__xnor2_2 _19972_ (.A(_03256_),
    .B(_03267_),
    .Y(_03278_));
 sky130_fd_sc_hd__and4_2 _19973_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[16]),
    .D(iX[17]),
    .X(_03289_));
 sky130_fd_sc_hd__a22oi_2 _19974_ (.A1(iY[4]),
    .A2(iX[16]),
    .B1(iX[17]),
    .B2(iY[3]),
    .Y(_03299_));
 sky130_fd_sc_hd__nor2_2 _19975_ (.A(_03289_),
    .B(_03299_),
    .Y(_03310_));
 sky130_fd_sc_hd__nand2_2 _19976_ (.A(iY[5]),
    .B(iX[15]),
    .Y(_03321_));
 sky130_fd_sc_hd__xnor2_2 _19977_ (.A(_03310_),
    .B(_03321_),
    .Y(_03332_));
 sky130_fd_sc_hd__xnor2_2 _19978_ (.A(_03278_),
    .B(_03332_),
    .Y(_03343_));
 sky130_fd_sc_hd__a21o_2 _19979_ (.A1(_03190_),
    .A2(_03201_),
    .B1(_03343_),
    .X(_03354_));
 sky130_fd_sc_hd__nand3_2 _19980_ (.A(_03190_),
    .B(_03201_),
    .C(_03343_),
    .Y(_03365_));
 sky130_fd_sc_hd__o21ba_2 _19981_ (.A1(_02500_),
    .A2(_02521_),
    .B1_N(_02489_),
    .X(_03376_));
 sky130_fd_sc_hd__o21ba_2 _19982_ (.A1(_02390_),
    .A2(_02412_),
    .B1_N(_02379_),
    .X(_03387_));
 sky130_fd_sc_hd__and4_2 _19983_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[13]),
    .D(iX[14]),
    .X(_03398_));
 sky130_fd_sc_hd__a22oi_2 _19984_ (.A1(iY[7]),
    .A2(iX[13]),
    .B1(iX[14]),
    .B2(iY[6]),
    .Y(_03409_));
 sky130_fd_sc_hd__nor2_2 _19985_ (.A(_03398_),
    .B(_03409_),
    .Y(_03420_));
 sky130_fd_sc_hd__nand2_2 _19986_ (.A(iY[8]),
    .B(iX[12]),
    .Y(_03431_));
 sky130_fd_sc_hd__xnor2_2 _19987_ (.A(_03420_),
    .B(_03431_),
    .Y(_03442_));
 sky130_fd_sc_hd__xnor2_2 _19988_ (.A(_03387_),
    .B(_03442_),
    .Y(_03453_));
 sky130_fd_sc_hd__xnor2_2 _19989_ (.A(_03376_),
    .B(_03453_),
    .Y(_03464_));
 sky130_fd_sc_hd__nand3_2 _19990_ (.A(_03354_),
    .B(_03365_),
    .C(_03464_),
    .Y(_03475_));
 sky130_fd_sc_hd__a21o_2 _19991_ (.A1(_03354_),
    .A2(_03365_),
    .B1(_03464_),
    .X(_03486_));
 sky130_fd_sc_hd__nand2_2 _19992_ (.A(_02445_),
    .B(_02565_),
    .Y(_03497_));
 sky130_fd_sc_hd__and3_2 _19993_ (.A(_03475_),
    .B(_03486_),
    .C(_03497_),
    .X(_03508_));
 sky130_fd_sc_hd__a21oi_2 _19994_ (.A1(_03475_),
    .A2(_03486_),
    .B1(_03497_),
    .Y(_03519_));
 sky130_fd_sc_hd__and2b_2 _19995_ (.A_N(_02181_),
    .B(_02170_),
    .X(_03530_));
 sky130_fd_sc_hd__or2b_2 _19996_ (.A(_02478_),
    .B_N(_02532_),
    .X(_03541_));
 sky130_fd_sc_hd__or2b_2 _19997_ (.A(_02467_),
    .B_N(_02543_),
    .X(_03552_));
 sky130_fd_sc_hd__and4_2 _19998_ (.A(iX[7]),
    .B(iX[8]),
    .C(iY[12]),
    .D(iY[13]),
    .X(_03563_));
 sky130_fd_sc_hd__a22oi_2 _19999_ (.A1(iX[8]),
    .A2(iY[12]),
    .B1(iY[13]),
    .B2(iX[7]),
    .Y(_03574_));
 sky130_fd_sc_hd__nor2_2 _20000_ (.A(_03563_),
    .B(_03574_),
    .Y(_03585_));
 sky130_fd_sc_hd__nand2_2 _20001_ (.A(iX[6]),
    .B(iY[14]),
    .Y(_03596_));
 sky130_fd_sc_hd__xnor2_2 _20002_ (.A(_03585_),
    .B(_03596_),
    .Y(_03607_));
 sky130_fd_sc_hd__and4_2 _20003_ (.A(iY[9]),
    .B(iX[10]),
    .C(iY[10]),
    .D(iX[11]),
    .X(_03618_));
 sky130_fd_sc_hd__a22oi_2 _20004_ (.A1(iX[10]),
    .A2(iY[10]),
    .B1(iX[11]),
    .B2(iY[9]),
    .Y(_03629_));
 sky130_fd_sc_hd__nor2_2 _20005_ (.A(_03618_),
    .B(_03629_),
    .Y(_03640_));
 sky130_fd_sc_hd__nand2_2 _20006_ (.A(iX[9]),
    .B(iY[11]),
    .Y(_03651_));
 sky130_fd_sc_hd__xnor2_2 _20007_ (.A(_03640_),
    .B(_03651_),
    .Y(_03662_));
 sky130_fd_sc_hd__o21ba_2 _20008_ (.A1(_02137_),
    .A2(_02159_),
    .B1_N(_02126_),
    .X(_03673_));
 sky130_fd_sc_hd__xnor2_2 _20009_ (.A(_03662_),
    .B(_03673_),
    .Y(_03684_));
 sky130_fd_sc_hd__and2_2 _20010_ (.A(_03607_),
    .B(_03684_),
    .X(_03694_));
 sky130_fd_sc_hd__nor2_2 _20011_ (.A(_03607_),
    .B(_03684_),
    .Y(_03705_));
 sky130_fd_sc_hd__or2_2 _20012_ (.A(_03694_),
    .B(_03705_),
    .X(_03716_));
 sky130_fd_sc_hd__a21o_2 _20013_ (.A1(_03541_),
    .A2(_03552_),
    .B1(_03716_),
    .X(_03727_));
 sky130_fd_sc_hd__nand3_2 _20014_ (.A(_03541_),
    .B(_03552_),
    .C(_03716_),
    .Y(_03738_));
 sky130_fd_sc_hd__o211ai_2 _20015_ (.A1(_03530_),
    .A2(_02203_),
    .B1(_03727_),
    .C1(_03738_),
    .Y(_03749_));
 sky130_fd_sc_hd__a211o_2 _20016_ (.A1(_03727_),
    .A2(_03738_),
    .B1(_03530_),
    .C1(_02203_),
    .X(_03760_));
 sky130_fd_sc_hd__a2bb2o_2 _20017_ (.A1_N(_03508_),
    .A2_N(_03519_),
    .B1(_03749_),
    .B2(_03760_),
    .X(_03771_));
 sky130_fd_sc_hd__or4bb_2 _20018_ (.A(_03508_),
    .B(_03519_),
    .C_N(_03749_),
    .D_N(_03760_),
    .X(_03782_));
 sky130_fd_sc_hd__o211a_2 _20019_ (.A1(_03179_),
    .A2(_02631_),
    .B1(_03771_),
    .C1(_03782_),
    .X(_03793_));
 sky130_fd_sc_hd__a211oi_2 _20020_ (.A1(_03771_),
    .A2(_03782_),
    .B1(_03179_),
    .C1(_02631_),
    .Y(_03804_));
 sky130_fd_sc_hd__and4_2 _20021_ (.A(iX[1]),
    .B(iX[2]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_03815_));
 sky130_fd_sc_hd__a22oi_2 _20022_ (.A1(iX[2]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[1]),
    .Y(_03826_));
 sky130_fd_sc_hd__nor2_2 _20023_ (.A(_03815_),
    .B(_03826_),
    .Y(_03837_));
 sky130_fd_sc_hd__nand2_2 _20024_ (.A(iX[0]),
    .B(iY[20]),
    .Y(_03848_));
 sky130_fd_sc_hd__xnor2_2 _20025_ (.A(_03837_),
    .B(_03848_),
    .Y(_03859_));
 sky130_fd_sc_hd__and2_2 _20026_ (.A(_02697_),
    .B(_03859_),
    .X(_03870_));
 sky130_fd_sc_hd__nor2_2 _20027_ (.A(_02697_),
    .B(_03859_),
    .Y(_03881_));
 sky130_fd_sc_hd__or2_2 _20028_ (.A(_03870_),
    .B(_03881_),
    .X(_03892_));
 sky130_fd_sc_hd__or2b_2 _20029_ (.A(_02730_),
    .B_N(_02785_),
    .X(_03903_));
 sky130_fd_sc_hd__a31o_2 _20030_ (.A1(iX[2]),
    .A2(iY[17]),
    .A3(_02763_),
    .B1(_02741_),
    .X(_03914_));
 sky130_fd_sc_hd__o21ba_2 _20031_ (.A1(_02083_),
    .A2(_02105_),
    .B1_N(_02072_),
    .X(_03925_));
 sky130_fd_sc_hd__and4_2 _20032_ (.A(iX[4]),
    .B(iX[5]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_03936_));
 sky130_fd_sc_hd__a22oi_2 _20033_ (.A1(iX[5]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[4]),
    .Y(_03947_));
 sky130_fd_sc_hd__nor2_2 _20034_ (.A(_03936_),
    .B(_03947_),
    .Y(_03958_));
 sky130_fd_sc_hd__nand2_2 _20035_ (.A(iX[3]),
    .B(iY[17]),
    .Y(_03969_));
 sky130_fd_sc_hd__xnor2_2 _20036_ (.A(_03958_),
    .B(_03969_),
    .Y(_03980_));
 sky130_fd_sc_hd__xnor2_2 _20037_ (.A(_03925_),
    .B(_03980_),
    .Y(_03991_));
 sky130_fd_sc_hd__xnor2_2 _20038_ (.A(_03914_),
    .B(_03991_),
    .Y(_04002_));
 sky130_fd_sc_hd__a21oi_2 _20039_ (.A1(_03903_),
    .A2(_02807_),
    .B1(_04002_),
    .Y(_04013_));
 sky130_fd_sc_hd__and3_2 _20040_ (.A(_03903_),
    .B(_02807_),
    .C(_04002_),
    .X(_04024_));
 sky130_fd_sc_hd__or3_2 _20041_ (.A(_03892_),
    .B(_04013_),
    .C(_04024_),
    .X(_04035_));
 sky130_fd_sc_hd__o21ai_2 _20042_ (.A1(_04013_),
    .A2(_04024_),
    .B1(_03892_),
    .Y(_04046_));
 sky130_fd_sc_hd__nand2_2 _20043_ (.A(_04035_),
    .B(_04046_),
    .Y(_04056_));
 sky130_fd_sc_hd__a21oi_2 _20044_ (.A1(_02236_),
    .A2(_02258_),
    .B1(_04056_),
    .Y(_04067_));
 sky130_fd_sc_hd__and3_2 _20045_ (.A(_02236_),
    .B(_02258_),
    .C(_04056_),
    .X(_04078_));
 sky130_fd_sc_hd__a211oi_2 _20046_ (.A1(_02840_),
    .A2(_02873_),
    .B1(_04067_),
    .C1(_04078_),
    .Y(_04089_));
 sky130_fd_sc_hd__o211a_2 _20047_ (.A1(_04067_),
    .A2(_04078_),
    .B1(_02840_),
    .C1(_02873_),
    .X(_04100_));
 sky130_fd_sc_hd__nor4_2 _20048_ (.A(_03793_),
    .B(_03804_),
    .C(_04089_),
    .D(_04100_),
    .Y(_04111_));
 sky130_fd_sc_hd__o22a_2 _20049_ (.A1(_03793_),
    .A2(_03804_),
    .B1(_04089_),
    .B2(_04100_),
    .X(_04122_));
 sky130_fd_sc_hd__a211oi_2 _20050_ (.A1(_02653_),
    .A2(_02949_),
    .B1(_04111_),
    .C1(_04122_),
    .Y(_04133_));
 sky130_fd_sc_hd__o211a_2 _20051_ (.A1(_04111_),
    .A2(_04122_),
    .B1(_02653_),
    .C1(_02949_),
    .X(_04144_));
 sky130_fd_sc_hd__and2b_2 _20052_ (.A_N(_02895_),
    .B(_02927_),
    .X(_04155_));
 sky130_fd_sc_hd__or3_2 _20053_ (.A(_04133_),
    .B(_04144_),
    .C(_04155_),
    .X(_04166_));
 sky130_fd_sc_hd__o21ai_2 _20054_ (.A1(_04133_),
    .A2(_04144_),
    .B1(_04155_),
    .Y(_04177_));
 sky130_fd_sc_hd__nand2_2 _20055_ (.A(_04166_),
    .B(_04177_),
    .Y(_04188_));
 sky130_fd_sc_hd__a21o_2 _20056_ (.A1(_02982_),
    .A2(_03026_),
    .B1(_02971_),
    .X(_04199_));
 sky130_fd_sc_hd__xnor2_2 _20057_ (.A(_04188_),
    .B(_04199_),
    .Y(_04210_));
 sky130_fd_sc_hd__nor3b_2 _20058_ (.A(_03037_),
    .B(_03048_),
    .C_N(_04210_),
    .Y(_04221_));
 sky130_fd_sc_hd__o21ba_2 _20059_ (.A1(_03037_),
    .A2(_03048_),
    .B1_N(_04210_),
    .X(_04232_));
 sky130_fd_sc_hd__and4bb_2 _20060_ (.A_N(_04221_),
    .B_N(_04232_),
    .C(_02017_),
    .D(_03059_),
    .X(_04243_));
 sky130_fd_sc_hd__o2bb2a_2 _20061_ (.A1_N(_02017_),
    .A2_N(_03059_),
    .B1(_04221_),
    .B2(_04232_),
    .X(_04254_));
 sky130_fd_sc_hd__nor2_2 _20062_ (.A(_04243_),
    .B(_04254_),
    .Y(_04265_));
 sky130_fd_sc_hd__nand2_2 _20063_ (.A(_03168_),
    .B(_04265_),
    .Y(_04276_));
 sky130_fd_sc_hd__or2_2 _20064_ (.A(_03168_),
    .B(_04265_),
    .X(_04287_));
 sky130_fd_sc_hd__and2_2 _20065_ (.A(_04276_),
    .B(_04287_),
    .X(_04298_));
 sky130_fd_sc_hd__buf_1 _20066_ (.A(_04298_),
    .X(oO[20]));
 sky130_fd_sc_hd__or2b_2 _20067_ (.A(_04188_),
    .B_N(_04199_),
    .X(_04319_));
 sky130_fd_sc_hd__and4bb_2 _20068_ (.A_N(_03508_),
    .B_N(_03519_),
    .C(_03749_),
    .D(_03760_),
    .X(_04330_));
 sky130_fd_sc_hd__or2b_2 _20069_ (.A(_03267_),
    .B_N(_03256_),
    .X(_04341_));
 sky130_fd_sc_hd__nand2_2 _20070_ (.A(_03278_),
    .B(_03332_),
    .Y(_04352_));
 sky130_fd_sc_hd__and4_2 _20071_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[20]),
    .D(iX[21]),
    .X(_04363_));
 sky130_fd_sc_hd__a22oi_2 _20072_ (.A1(iY[1]),
    .A2(iX[20]),
    .B1(iX[21]),
    .B2(iY[0]),
    .Y(_04374_));
 sky130_fd_sc_hd__nor2_2 _20073_ (.A(_04363_),
    .B(_04374_),
    .Y(_04385_));
 sky130_fd_sc_hd__nand2_2 _20074_ (.A(iY[2]),
    .B(iX[19]),
    .Y(_04396_));
 sky130_fd_sc_hd__xnor2_2 _20075_ (.A(_04385_),
    .B(_04396_),
    .Y(_04407_));
 sky130_fd_sc_hd__o21ba_2 _20076_ (.A1(_03223_),
    .A2(_03245_),
    .B1_N(_03212_),
    .X(_04418_));
 sky130_fd_sc_hd__xnor2_2 _20077_ (.A(_04407_),
    .B(_04418_),
    .Y(_04429_));
 sky130_fd_sc_hd__and4_2 _20078_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[17]),
    .D(iX[18]),
    .X(_04439_));
 sky130_fd_sc_hd__a22oi_2 _20079_ (.A1(iY[4]),
    .A2(iX[17]),
    .B1(iX[18]),
    .B2(iY[3]),
    .Y(_04450_));
 sky130_fd_sc_hd__nor2_2 _20080_ (.A(_04439_),
    .B(_04450_),
    .Y(_04461_));
 sky130_fd_sc_hd__nand2_2 _20081_ (.A(iY[5]),
    .B(iX[16]),
    .Y(_04472_));
 sky130_fd_sc_hd__xnor2_2 _20082_ (.A(_04461_),
    .B(_04472_),
    .Y(_04483_));
 sky130_fd_sc_hd__xnor2_2 _20083_ (.A(_04429_),
    .B(_04483_),
    .Y(_04494_));
 sky130_fd_sc_hd__a21o_2 _20084_ (.A1(_04341_),
    .A2(_04352_),
    .B1(_04494_),
    .X(_04505_));
 sky130_fd_sc_hd__nand3_2 _20085_ (.A(_04341_),
    .B(_04352_),
    .C(_04494_),
    .Y(_04516_));
 sky130_fd_sc_hd__o21ba_2 _20086_ (.A1(_03409_),
    .A2(_03431_),
    .B1_N(_03398_),
    .X(_04527_));
 sky130_fd_sc_hd__o21ba_2 _20087_ (.A1(_03299_),
    .A2(_03321_),
    .B1_N(_03289_),
    .X(_04538_));
 sky130_fd_sc_hd__and4_2 _20088_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[14]),
    .D(iX[15]),
    .X(_04549_));
 sky130_fd_sc_hd__a22oi_2 _20089_ (.A1(iY[7]),
    .A2(iX[14]),
    .B1(iX[15]),
    .B2(iY[6]),
    .Y(_04560_));
 sky130_fd_sc_hd__nor2_2 _20090_ (.A(_04549_),
    .B(_04560_),
    .Y(_04571_));
 sky130_fd_sc_hd__nand2_2 _20091_ (.A(iY[8]),
    .B(iX[13]),
    .Y(_04582_));
 sky130_fd_sc_hd__xnor2_2 _20092_ (.A(_04571_),
    .B(_04582_),
    .Y(_04593_));
 sky130_fd_sc_hd__xnor2_2 _20093_ (.A(_04538_),
    .B(_04593_),
    .Y(_04604_));
 sky130_fd_sc_hd__xnor2_2 _20094_ (.A(_04527_),
    .B(_04604_),
    .Y(_04615_));
 sky130_fd_sc_hd__nand3_2 _20095_ (.A(_04505_),
    .B(_04516_),
    .C(_04615_),
    .Y(_04626_));
 sky130_fd_sc_hd__a21o_2 _20096_ (.A1(_04505_),
    .A2(_04516_),
    .B1(_04615_),
    .X(_04637_));
 sky130_fd_sc_hd__nand2_2 _20097_ (.A(_03354_),
    .B(_03475_),
    .Y(_04648_));
 sky130_fd_sc_hd__and3_2 _20098_ (.A(_04626_),
    .B(_04637_),
    .C(_04648_),
    .X(_04659_));
 sky130_fd_sc_hd__a21oi_2 _20099_ (.A1(_04626_),
    .A2(_04637_),
    .B1(_04648_),
    .Y(_04670_));
 sky130_fd_sc_hd__and2b_2 _20100_ (.A_N(_03673_),
    .B(_03662_),
    .X(_04681_));
 sky130_fd_sc_hd__or2b_2 _20101_ (.A(_03387_),
    .B_N(_03442_),
    .X(_04692_));
 sky130_fd_sc_hd__or2b_2 _20102_ (.A(_03376_),
    .B_N(_03453_),
    .X(_04703_));
 sky130_fd_sc_hd__and4_2 _20103_ (.A(iX[8]),
    .B(iX[9]),
    .C(iY[12]),
    .D(iY[13]),
    .X(_04714_));
 sky130_fd_sc_hd__a22oi_2 _20104_ (.A1(iX[9]),
    .A2(iY[12]),
    .B1(iY[13]),
    .B2(iX[8]),
    .Y(_04725_));
 sky130_fd_sc_hd__nor2_2 _20105_ (.A(_04714_),
    .B(_04725_),
    .Y(_04736_));
 sky130_fd_sc_hd__nand2_2 _20106_ (.A(iX[7]),
    .B(iY[14]),
    .Y(_04747_));
 sky130_fd_sc_hd__xnor2_2 _20107_ (.A(_04736_),
    .B(_04747_),
    .Y(_04758_));
 sky130_fd_sc_hd__and4_2 _20108_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[11]),
    .D(iX[12]),
    .X(_04768_));
 sky130_fd_sc_hd__a22oi_2 _20109_ (.A1(iY[10]),
    .A2(iX[11]),
    .B1(iX[12]),
    .B2(iY[9]),
    .Y(_04779_));
 sky130_fd_sc_hd__nor2_2 _20110_ (.A(_04768_),
    .B(_04779_),
    .Y(_04790_));
 sky130_fd_sc_hd__nand2_2 _20111_ (.A(iX[10]),
    .B(iY[11]),
    .Y(_04801_));
 sky130_fd_sc_hd__xnor2_2 _20112_ (.A(_04790_),
    .B(_04801_),
    .Y(_04812_));
 sky130_fd_sc_hd__o21ba_2 _20113_ (.A1(_03629_),
    .A2(_03651_),
    .B1_N(_03618_),
    .X(_04823_));
 sky130_fd_sc_hd__xnor2_2 _20114_ (.A(_04812_),
    .B(_04823_),
    .Y(_04834_));
 sky130_fd_sc_hd__and2_2 _20115_ (.A(_04758_),
    .B(_04834_),
    .X(_04845_));
 sky130_fd_sc_hd__nor2_2 _20116_ (.A(_04758_),
    .B(_04834_),
    .Y(_04856_));
 sky130_fd_sc_hd__or2_2 _20117_ (.A(_04845_),
    .B(_04856_),
    .X(_04867_));
 sky130_fd_sc_hd__a21o_2 _20118_ (.A1(_04692_),
    .A2(_04703_),
    .B1(_04867_),
    .X(_04878_));
 sky130_fd_sc_hd__nand3_2 _20119_ (.A(_04692_),
    .B(_04703_),
    .C(_04867_),
    .Y(_04889_));
 sky130_fd_sc_hd__o211ai_2 _20120_ (.A1(_04681_),
    .A2(_03694_),
    .B1(_04878_),
    .C1(_04889_),
    .Y(_04900_));
 sky130_fd_sc_hd__a211o_2 _20121_ (.A1(_04878_),
    .A2(_04889_),
    .B1(_04681_),
    .C1(_03694_),
    .X(_04911_));
 sky130_fd_sc_hd__a2bb2o_2 _20122_ (.A1_N(_04659_),
    .A2_N(_04670_),
    .B1(_04900_),
    .B2(_04911_),
    .X(_04922_));
 sky130_fd_sc_hd__or4bb_2 _20123_ (.A(_04659_),
    .B(_04670_),
    .C_N(_04900_),
    .D_N(_04911_),
    .X(_04933_));
 sky130_fd_sc_hd__o211ai_2 _20124_ (.A1(_03508_),
    .A2(_04330_),
    .B1(_04922_),
    .C1(_04933_),
    .Y(_04944_));
 sky130_fd_sc_hd__a211o_2 _20125_ (.A1(_04922_),
    .A2(_04933_),
    .B1(_03508_),
    .C1(_04330_),
    .X(_04955_));
 sky130_fd_sc_hd__inv_2 _20126_ (.A(_04013_),
    .Y(_04966_));
 sky130_fd_sc_hd__and4_2 _20127_ (.A(iX[2]),
    .B(iX[3]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_04977_));
 sky130_fd_sc_hd__a22oi_2 _20128_ (.A1(iX[3]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[2]),
    .Y(_04988_));
 sky130_fd_sc_hd__nor2_2 _20129_ (.A(_04977_),
    .B(_04988_),
    .Y(_04999_));
 sky130_fd_sc_hd__nand2_2 _20130_ (.A(iX[1]),
    .B(iY[20]),
    .Y(_05010_));
 sky130_fd_sc_hd__xnor2_2 _20131_ (.A(_04999_),
    .B(_05010_),
    .Y(_05021_));
 sky130_fd_sc_hd__o21ba_2 _20132_ (.A1(_03826_),
    .A2(_03848_),
    .B1_N(_03815_),
    .X(_05032_));
 sky130_fd_sc_hd__xnor2_2 _20133_ (.A(_05021_),
    .B(_05032_),
    .Y(_05043_));
 sky130_fd_sc_hd__nand2_2 _20134_ (.A(iX[0]),
    .B(iY[21]),
    .Y(_05054_));
 sky130_fd_sc_hd__xor2_2 _20135_ (.A(_05043_),
    .B(_05054_),
    .X(_05065_));
 sky130_fd_sc_hd__or2b_2 _20136_ (.A(_03925_),
    .B_N(_03980_),
    .X(_05076_));
 sky130_fd_sc_hd__nand2_2 _20137_ (.A(_03914_),
    .B(_03991_),
    .Y(_05087_));
 sky130_fd_sc_hd__a31o_2 _20138_ (.A1(iX[3]),
    .A2(iY[17]),
    .A3(_03958_),
    .B1(_03936_),
    .X(_05098_));
 sky130_fd_sc_hd__o21ba_2 _20139_ (.A1(_03574_),
    .A2(_03596_),
    .B1_N(_03563_),
    .X(_05108_));
 sky130_fd_sc_hd__and4_2 _20140_ (.A(iX[5]),
    .B(iX[6]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_05119_));
 sky130_fd_sc_hd__a22oi_2 _20141_ (.A1(iX[6]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[5]),
    .Y(_05130_));
 sky130_fd_sc_hd__nor2_2 _20142_ (.A(_05119_),
    .B(_05130_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand2_2 _20143_ (.A(iX[4]),
    .B(iY[17]),
    .Y(_05152_));
 sky130_fd_sc_hd__xnor2_2 _20144_ (.A(_05141_),
    .B(_05152_),
    .Y(_05163_));
 sky130_fd_sc_hd__xnor2_2 _20145_ (.A(_05108_),
    .B(_05163_),
    .Y(_05174_));
 sky130_fd_sc_hd__xnor2_2 _20146_ (.A(_05098_),
    .B(_05174_),
    .Y(_05185_));
 sky130_fd_sc_hd__a21oi_2 _20147_ (.A1(_05076_),
    .A2(_05087_),
    .B1(_05185_),
    .Y(_05196_));
 sky130_fd_sc_hd__and3_2 _20148_ (.A(_05076_),
    .B(_05087_),
    .C(_05185_),
    .X(_05207_));
 sky130_fd_sc_hd__or3_2 _20149_ (.A(_05065_),
    .B(_05196_),
    .C(_05207_),
    .X(_05218_));
 sky130_fd_sc_hd__o21ai_2 _20150_ (.A1(_05196_),
    .A2(_05207_),
    .B1(_05065_),
    .Y(_05229_));
 sky130_fd_sc_hd__nand2_2 _20151_ (.A(_05218_),
    .B(_05229_),
    .Y(_05240_));
 sky130_fd_sc_hd__a21oi_2 _20152_ (.A1(_03727_),
    .A2(_03749_),
    .B1(_05240_),
    .Y(_05251_));
 sky130_fd_sc_hd__and3_2 _20153_ (.A(_03727_),
    .B(_03749_),
    .C(_05240_),
    .X(_05262_));
 sky130_fd_sc_hd__a211oi_2 _20154_ (.A1(_04966_),
    .A2(_04035_),
    .B1(_05251_),
    .C1(_05262_),
    .Y(_05273_));
 sky130_fd_sc_hd__o211a_2 _20155_ (.A1(_05251_),
    .A2(_05262_),
    .B1(_04966_),
    .C1(_04035_),
    .X(_05284_));
 sky130_fd_sc_hd__nor2_2 _20156_ (.A(_05273_),
    .B(_05284_),
    .Y(_05295_));
 sky130_fd_sc_hd__nand3_2 _20157_ (.A(_04944_),
    .B(_04955_),
    .C(_05295_),
    .Y(_05306_));
 sky130_fd_sc_hd__a21o_2 _20158_ (.A1(_04944_),
    .A2(_04955_),
    .B1(_05295_),
    .X(_05317_));
 sky130_fd_sc_hd__o211ai_2 _20159_ (.A1(_03793_),
    .A2(_04111_),
    .B1(_05306_),
    .C1(_05317_),
    .Y(_05328_));
 sky130_fd_sc_hd__a211o_2 _20160_ (.A1(_05306_),
    .A2(_05317_),
    .B1(_03793_),
    .C1(_04111_),
    .X(_05339_));
 sky130_fd_sc_hd__o21ai_2 _20161_ (.A1(_04067_),
    .A2(_04089_),
    .B1(_03870_),
    .Y(_05350_));
 sky130_fd_sc_hd__or3_2 _20162_ (.A(_03870_),
    .B(_04067_),
    .C(_04089_),
    .X(_05361_));
 sky130_fd_sc_hd__and2_2 _20163_ (.A(_05350_),
    .B(_05361_),
    .X(_05372_));
 sky130_fd_sc_hd__nand3_2 _20164_ (.A(_05328_),
    .B(_05339_),
    .C(_05372_),
    .Y(_05383_));
 sky130_fd_sc_hd__a21o_2 _20165_ (.A1(_05328_),
    .A2(_05339_),
    .B1(_05372_),
    .X(_05394_));
 sky130_fd_sc_hd__nand2_2 _20166_ (.A(_05383_),
    .B(_05394_),
    .Y(_05405_));
 sky130_fd_sc_hd__o21ba_2 _20167_ (.A1(_04144_),
    .A2(_04155_),
    .B1_N(_04133_),
    .X(_05416_));
 sky130_fd_sc_hd__xnor2_2 _20168_ (.A(_05405_),
    .B(_05416_),
    .Y(_05426_));
 sky130_fd_sc_hd__xor2_2 _20169_ (.A(_04319_),
    .B(_05426_),
    .X(_05437_));
 sky130_fd_sc_hd__and2_2 _20170_ (.A(_04221_),
    .B(_05437_),
    .X(_05448_));
 sky130_fd_sc_hd__nor2_2 _20171_ (.A(_04221_),
    .B(_05437_),
    .Y(_05459_));
 sky130_fd_sc_hd__or2_2 _20172_ (.A(_05448_),
    .B(_05459_),
    .X(_05470_));
 sky130_fd_sc_hd__and3b_2 _20173_ (.A_N(_04243_),
    .B(_04276_),
    .C(_05470_),
    .X(_05481_));
 sky130_fd_sc_hd__and2_2 _20174_ (.A(_04243_),
    .B(_05437_),
    .X(_05492_));
 sky130_fd_sc_hd__o21bai_2 _20175_ (.A1(_04276_),
    .A2(_05470_),
    .B1_N(_05492_),
    .Y(_05503_));
 sky130_fd_sc_hd__nor2_2 _20176_ (.A(_05481_),
    .B(_05503_),
    .Y(oO[21]));
 sky130_fd_sc_hd__nor2_2 _20177_ (.A(_04319_),
    .B(_05426_),
    .Y(_05524_));
 sky130_fd_sc_hd__or2_2 _20178_ (.A(_05405_),
    .B(_05416_),
    .X(_05535_));
 sky130_fd_sc_hd__and4bb_2 _20179_ (.A_N(_04659_),
    .B_N(_04670_),
    .C(_04900_),
    .D(_04911_),
    .X(_05546_));
 sky130_fd_sc_hd__or2b_2 _20180_ (.A(_04418_),
    .B_N(_04407_),
    .X(_05557_));
 sky130_fd_sc_hd__nand2_2 _20181_ (.A(_04429_),
    .B(_04483_),
    .Y(_05568_));
 sky130_fd_sc_hd__and4_2 _20182_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[21]),
    .D(iX[22]),
    .X(_05579_));
 sky130_fd_sc_hd__a22oi_2 _20183_ (.A1(iY[1]),
    .A2(iX[21]),
    .B1(iX[22]),
    .B2(iY[0]),
    .Y(_05590_));
 sky130_fd_sc_hd__nor2_2 _20184_ (.A(_05579_),
    .B(_05590_),
    .Y(_05601_));
 sky130_fd_sc_hd__nand2_2 _20185_ (.A(iY[2]),
    .B(iX[20]),
    .Y(_05612_));
 sky130_fd_sc_hd__xnor2_2 _20186_ (.A(_05601_),
    .B(_05612_),
    .Y(_05623_));
 sky130_fd_sc_hd__o21ba_2 _20187_ (.A1(_04374_),
    .A2(_04396_),
    .B1_N(_04363_),
    .X(_05634_));
 sky130_fd_sc_hd__xnor2_2 _20188_ (.A(_05623_),
    .B(_05634_),
    .Y(_05645_));
 sky130_fd_sc_hd__and4_2 _20189_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[18]),
    .D(iX[19]),
    .X(_05656_));
 sky130_fd_sc_hd__a22oi_2 _20190_ (.A1(iY[4]),
    .A2(iX[18]),
    .B1(iX[19]),
    .B2(iY[3]),
    .Y(_05667_));
 sky130_fd_sc_hd__nor2_2 _20191_ (.A(_05656_),
    .B(_05667_),
    .Y(_05678_));
 sky130_fd_sc_hd__nand2_2 _20192_ (.A(iY[5]),
    .B(iX[17]),
    .Y(_05689_));
 sky130_fd_sc_hd__xnor2_2 _20193_ (.A(_05678_),
    .B(_05689_),
    .Y(_05700_));
 sky130_fd_sc_hd__xnor2_2 _20194_ (.A(_05645_),
    .B(_05700_),
    .Y(_05711_));
 sky130_fd_sc_hd__a21o_2 _20195_ (.A1(_05557_),
    .A2(_05568_),
    .B1(_05711_),
    .X(_05722_));
 sky130_fd_sc_hd__nand3_2 _20196_ (.A(_05557_),
    .B(_05568_),
    .C(_05711_),
    .Y(_05733_));
 sky130_fd_sc_hd__o21ba_2 _20197_ (.A1(_04560_),
    .A2(_04582_),
    .B1_N(_04549_),
    .X(_05744_));
 sky130_fd_sc_hd__o21ba_2 _20198_ (.A1(_04450_),
    .A2(_04472_),
    .B1_N(_04439_),
    .X(_05755_));
 sky130_fd_sc_hd__and4_2 _20199_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[15]),
    .D(iX[16]),
    .X(_05766_));
 sky130_fd_sc_hd__a22oi_2 _20200_ (.A1(iY[7]),
    .A2(iX[15]),
    .B1(iX[16]),
    .B2(iY[6]),
    .Y(_05777_));
 sky130_fd_sc_hd__nor2_2 _20201_ (.A(_05766_),
    .B(_05777_),
    .Y(_05787_));
 sky130_fd_sc_hd__nand2_2 _20202_ (.A(iY[8]),
    .B(iX[14]),
    .Y(_05798_));
 sky130_fd_sc_hd__xnor2_2 _20203_ (.A(_05787_),
    .B(_05798_),
    .Y(_05809_));
 sky130_fd_sc_hd__xnor2_2 _20204_ (.A(_05755_),
    .B(_05809_),
    .Y(_05820_));
 sky130_fd_sc_hd__xnor2_2 _20205_ (.A(_05744_),
    .B(_05820_),
    .Y(_05831_));
 sky130_fd_sc_hd__nand3_2 _20206_ (.A(_05722_),
    .B(_05733_),
    .C(_05831_),
    .Y(_05842_));
 sky130_fd_sc_hd__a21o_2 _20207_ (.A1(_05722_),
    .A2(_05733_),
    .B1(_05831_),
    .X(_05853_));
 sky130_fd_sc_hd__nand2_2 _20208_ (.A(_04505_),
    .B(_04626_),
    .Y(_05864_));
 sky130_fd_sc_hd__and3_2 _20209_ (.A(_05842_),
    .B(_05853_),
    .C(_05864_),
    .X(_05875_));
 sky130_fd_sc_hd__a21oi_2 _20210_ (.A1(_05842_),
    .A2(_05853_),
    .B1(_05864_),
    .Y(_05886_));
 sky130_fd_sc_hd__and2b_2 _20211_ (.A_N(_04823_),
    .B(_04812_),
    .X(_05897_));
 sky130_fd_sc_hd__or2b_2 _20212_ (.A(_04538_),
    .B_N(_04593_),
    .X(_05908_));
 sky130_fd_sc_hd__or2b_2 _20213_ (.A(_04527_),
    .B_N(_04604_),
    .X(_05919_));
 sky130_fd_sc_hd__and4_2 _20214_ (.A(iX[9]),
    .B(iX[10]),
    .C(iY[12]),
    .D(iY[13]),
    .X(_05930_));
 sky130_fd_sc_hd__a22oi_2 _20215_ (.A1(iX[10]),
    .A2(iY[12]),
    .B1(iY[13]),
    .B2(iX[9]),
    .Y(_05941_));
 sky130_fd_sc_hd__nor2_2 _20216_ (.A(_05930_),
    .B(_05941_),
    .Y(_05952_));
 sky130_fd_sc_hd__nand2_2 _20217_ (.A(iX[8]),
    .B(iY[14]),
    .Y(_05963_));
 sky130_fd_sc_hd__xnor2_2 _20218_ (.A(_05952_),
    .B(_05963_),
    .Y(_05974_));
 sky130_fd_sc_hd__and4_2 _20219_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[12]),
    .D(iX[13]),
    .X(_05985_));
 sky130_fd_sc_hd__a22oi_2 _20220_ (.A1(iY[10]),
    .A2(iX[12]),
    .B1(iX[13]),
    .B2(iY[9]),
    .Y(_05996_));
 sky130_fd_sc_hd__nor2_2 _20221_ (.A(_05985_),
    .B(_05996_),
    .Y(_06007_));
 sky130_fd_sc_hd__nand2_2 _20222_ (.A(iX[11]),
    .B(iY[11]),
    .Y(_06018_));
 sky130_fd_sc_hd__xnor2_2 _20223_ (.A(_06007_),
    .B(_06018_),
    .Y(_06029_));
 sky130_fd_sc_hd__o21ba_2 _20224_ (.A1(_04779_),
    .A2(_04801_),
    .B1_N(_04768_),
    .X(_06040_));
 sky130_fd_sc_hd__xnor2_2 _20225_ (.A(_06029_),
    .B(_06040_),
    .Y(_06051_));
 sky130_fd_sc_hd__and2_2 _20226_ (.A(_05974_),
    .B(_06051_),
    .X(_06062_));
 sky130_fd_sc_hd__nor2_2 _20227_ (.A(_05974_),
    .B(_06051_),
    .Y(_06073_));
 sky130_fd_sc_hd__or2_2 _20228_ (.A(_06062_),
    .B(_06073_),
    .X(_06083_));
 sky130_fd_sc_hd__a21o_2 _20229_ (.A1(_05908_),
    .A2(_05919_),
    .B1(_06083_),
    .X(_06094_));
 sky130_fd_sc_hd__nand3_2 _20230_ (.A(_05908_),
    .B(_05919_),
    .C(_06083_),
    .Y(_06105_));
 sky130_fd_sc_hd__o211ai_2 _20231_ (.A1(_05897_),
    .A2(_04845_),
    .B1(_06094_),
    .C1(_06105_),
    .Y(_06116_));
 sky130_fd_sc_hd__a211o_2 _20232_ (.A1(_06094_),
    .A2(_06105_),
    .B1(_05897_),
    .C1(_04845_),
    .X(_06127_));
 sky130_fd_sc_hd__a2bb2o_2 _20233_ (.A1_N(_05875_),
    .A2_N(_05886_),
    .B1(_06116_),
    .B2(_06127_),
    .X(_06138_));
 sky130_fd_sc_hd__or4bb_2 _20234_ (.A(_05875_),
    .B(_05886_),
    .C_N(_06116_),
    .D_N(_06127_),
    .X(_06149_));
 sky130_fd_sc_hd__o211a_2 _20235_ (.A1(_04659_),
    .A2(_05546_),
    .B1(_06138_),
    .C1(_06149_),
    .X(_06160_));
 sky130_fd_sc_hd__a211oi_2 _20236_ (.A1(_06138_),
    .A2(_06149_),
    .B1(_04659_),
    .C1(_05546_),
    .Y(_06171_));
 sky130_fd_sc_hd__and2b_2 _20237_ (.A_N(_05196_),
    .B(_05218_),
    .X(_06182_));
 sky130_fd_sc_hd__a22oi_2 _20238_ (.A1(iX[1]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[0]),
    .Y(_06193_));
 sky130_fd_sc_hd__and4_2 _20239_ (.A(iX[0]),
    .B(iX[1]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_06204_));
 sky130_fd_sc_hd__or2_2 _20240_ (.A(_06193_),
    .B(_06204_),
    .X(_06215_));
 sky130_fd_sc_hd__and4_2 _20241_ (.A(iX[3]),
    .B(iX[4]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_06226_));
 sky130_fd_sc_hd__a22o_2 _20242_ (.A1(iX[4]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[3]),
    .X(_06237_));
 sky130_fd_sc_hd__and2b_2 _20243_ (.A_N(_06226_),
    .B(_06237_),
    .X(_06248_));
 sky130_fd_sc_hd__nand2_2 _20244_ (.A(iX[2]),
    .B(iY[20]),
    .Y(_06259_));
 sky130_fd_sc_hd__xnor2_2 _20245_ (.A(_06248_),
    .B(_06259_),
    .Y(_06270_));
 sky130_fd_sc_hd__o21ba_2 _20246_ (.A1(_04988_),
    .A2(_05010_),
    .B1_N(_04977_),
    .X(_06281_));
 sky130_fd_sc_hd__xnor2_2 _20247_ (.A(_06270_),
    .B(_06281_),
    .Y(_06292_));
 sky130_fd_sc_hd__xnor2_2 _20248_ (.A(_06215_),
    .B(_06292_),
    .Y(_06303_));
 sky130_fd_sc_hd__or2b_2 _20249_ (.A(_05108_),
    .B_N(_05163_),
    .X(_06314_));
 sky130_fd_sc_hd__nand2_2 _20250_ (.A(_05098_),
    .B(_05174_),
    .Y(_06325_));
 sky130_fd_sc_hd__a31o_2 _20251_ (.A1(iX[4]),
    .A2(iY[17]),
    .A3(_05141_),
    .B1(_05119_),
    .X(_06336_));
 sky130_fd_sc_hd__o21ba_2 _20252_ (.A1(_04725_),
    .A2(_04747_),
    .B1_N(_04714_),
    .X(_06347_));
 sky130_fd_sc_hd__and4_2 _20253_ (.A(iX[6]),
    .B(iX[7]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_06358_));
 sky130_fd_sc_hd__a22oi_2 _20254_ (.A1(iX[7]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[6]),
    .Y(_06369_));
 sky130_fd_sc_hd__nor2_2 _20255_ (.A(_06358_),
    .B(_06369_),
    .Y(_06379_));
 sky130_fd_sc_hd__nand2_2 _20256_ (.A(iX[5]),
    .B(iY[17]),
    .Y(_06390_));
 sky130_fd_sc_hd__xnor2_2 _20257_ (.A(_06379_),
    .B(_06390_),
    .Y(_06401_));
 sky130_fd_sc_hd__xnor2_2 _20258_ (.A(_06347_),
    .B(_06401_),
    .Y(_06412_));
 sky130_fd_sc_hd__xnor2_2 _20259_ (.A(_06336_),
    .B(_06412_),
    .Y(_06423_));
 sky130_fd_sc_hd__a21o_2 _20260_ (.A1(_06314_),
    .A2(_06325_),
    .B1(_06423_),
    .X(_06434_));
 sky130_fd_sc_hd__nand3_2 _20261_ (.A(_06314_),
    .B(_06325_),
    .C(_06423_),
    .Y(_06445_));
 sky130_fd_sc_hd__and3_2 _20262_ (.A(_06303_),
    .B(_06434_),
    .C(_06445_),
    .X(_06456_));
 sky130_fd_sc_hd__a21oi_2 _20263_ (.A1(_06434_),
    .A2(_06445_),
    .B1(_06303_),
    .Y(_06467_));
 sky130_fd_sc_hd__a211o_2 _20264_ (.A1(_04878_),
    .A2(_04900_),
    .B1(_06456_),
    .C1(_06467_),
    .X(_06478_));
 sky130_fd_sc_hd__o211ai_2 _20265_ (.A1(_06456_),
    .A2(_06467_),
    .B1(_04878_),
    .C1(_04900_),
    .Y(_06489_));
 sky130_fd_sc_hd__nand2_2 _20266_ (.A(_06478_),
    .B(_06489_),
    .Y(_06500_));
 sky130_fd_sc_hd__xor2_2 _20267_ (.A(_06182_),
    .B(_06500_),
    .X(_06511_));
 sky130_fd_sc_hd__nor3b_2 _20268_ (.A(_06160_),
    .B(_06171_),
    .C_N(_06511_),
    .Y(_06522_));
 sky130_fd_sc_hd__o21ba_2 _20269_ (.A1(_06160_),
    .A2(_06171_),
    .B1_N(_06511_),
    .X(_06533_));
 sky130_fd_sc_hd__a211o_2 _20270_ (.A1(_04944_),
    .A2(_05306_),
    .B1(_06522_),
    .C1(_06533_),
    .X(_06544_));
 sky130_fd_sc_hd__o211ai_2 _20271_ (.A1(_06522_),
    .A2(_06533_),
    .B1(_04944_),
    .C1(_05306_),
    .Y(_06555_));
 sky130_fd_sc_hd__and2b_2 _20272_ (.A_N(_05032_),
    .B(_05021_),
    .X(_06566_));
 sky130_fd_sc_hd__a31oi_2 _20273_ (.A1(iX[0]),
    .A2(iY[21]),
    .A3(_05043_),
    .B1(_06566_),
    .Y(_06577_));
 sky130_fd_sc_hd__o21ba_2 _20274_ (.A1(_05251_),
    .A2(_05273_),
    .B1_N(_06577_),
    .X(_06588_));
 sky130_fd_sc_hd__or3b_2 _20275_ (.A(_05251_),
    .B(_05273_),
    .C_N(_06577_),
    .X(_06599_));
 sky130_fd_sc_hd__and2b_2 _20276_ (.A_N(_06588_),
    .B(_06599_),
    .X(_06610_));
 sky130_fd_sc_hd__and3_2 _20277_ (.A(_06544_),
    .B(_06555_),
    .C(_06610_),
    .X(_06621_));
 sky130_fd_sc_hd__a21oi_2 _20278_ (.A1(_06544_),
    .A2(_06555_),
    .B1(_06610_),
    .Y(_06632_));
 sky130_fd_sc_hd__nor2_2 _20279_ (.A(_06621_),
    .B(_06632_),
    .Y(_06643_));
 sky130_fd_sc_hd__nand2_2 _20280_ (.A(_05328_),
    .B(_05383_),
    .Y(_06654_));
 sky130_fd_sc_hd__xnor2_2 _20281_ (.A(_06643_),
    .B(_06654_),
    .Y(_06664_));
 sky130_fd_sc_hd__xnor2_2 _20282_ (.A(_05350_),
    .B(_06664_),
    .Y(_06675_));
 sky130_fd_sc_hd__xor2_2 _20283_ (.A(_05535_),
    .B(_06675_),
    .X(_06686_));
 sky130_fd_sc_hd__and2_2 _20284_ (.A(_05524_),
    .B(_06686_),
    .X(_06697_));
 sky130_fd_sc_hd__nor2_2 _20285_ (.A(_05524_),
    .B(_06686_),
    .Y(_06708_));
 sky130_fd_sc_hd__nor2_2 _20286_ (.A(_06697_),
    .B(_06708_),
    .Y(_06719_));
 sky130_fd_sc_hd__nor2_2 _20287_ (.A(_05448_),
    .B(_05503_),
    .Y(_06730_));
 sky130_fd_sc_hd__xnor2_2 _20288_ (.A(_06719_),
    .B(_06730_),
    .Y(oO[22]));
 sky130_fd_sc_hd__nor2_2 _20289_ (.A(_05535_),
    .B(_06675_),
    .Y(_06751_));
 sky130_fd_sc_hd__inv_2 _20290_ (.A(_06621_),
    .Y(_06762_));
 sky130_fd_sc_hd__inv_2 _20291_ (.A(_05875_),
    .Y(_06773_));
 sky130_fd_sc_hd__or2b_2 _20292_ (.A(_05634_),
    .B_N(_05623_),
    .X(_06784_));
 sky130_fd_sc_hd__nand2_2 _20293_ (.A(_05645_),
    .B(_05700_),
    .Y(_06795_));
 sky130_fd_sc_hd__and4_2 _20294_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[22]),
    .D(iX[23]),
    .X(_06806_));
 sky130_fd_sc_hd__a22oi_2 _20295_ (.A1(iY[1]),
    .A2(iX[22]),
    .B1(iX[23]),
    .B2(iY[0]),
    .Y(_06817_));
 sky130_fd_sc_hd__nor2_2 _20296_ (.A(_06806_),
    .B(_06817_),
    .Y(_06828_));
 sky130_fd_sc_hd__nand2_2 _20297_ (.A(iY[2]),
    .B(iX[21]),
    .Y(_06839_));
 sky130_fd_sc_hd__xnor2_2 _20298_ (.A(_06828_),
    .B(_06839_),
    .Y(_06850_));
 sky130_fd_sc_hd__o21ba_2 _20299_ (.A1(_05590_),
    .A2(_05612_),
    .B1_N(_05579_),
    .X(_06861_));
 sky130_fd_sc_hd__xnor2_2 _20300_ (.A(_06850_),
    .B(_06861_),
    .Y(_06872_));
 sky130_fd_sc_hd__and4_2 _20301_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[19]),
    .D(iX[20]),
    .X(_06883_));
 sky130_fd_sc_hd__a22oi_2 _20302_ (.A1(iY[4]),
    .A2(iX[19]),
    .B1(iX[20]),
    .B2(iY[3]),
    .Y(_06894_));
 sky130_fd_sc_hd__nor2_2 _20303_ (.A(_06883_),
    .B(_06894_),
    .Y(_06905_));
 sky130_fd_sc_hd__nand2_2 _20304_ (.A(iY[5]),
    .B(iX[18]),
    .Y(_06916_));
 sky130_fd_sc_hd__xnor2_2 _20305_ (.A(_06905_),
    .B(_06916_),
    .Y(_06927_));
 sky130_fd_sc_hd__xnor2_2 _20306_ (.A(_06872_),
    .B(_06927_),
    .Y(_06938_));
 sky130_fd_sc_hd__a21o_2 _20307_ (.A1(_06784_),
    .A2(_06795_),
    .B1(_06938_),
    .X(_06948_));
 sky130_fd_sc_hd__nand3_2 _20308_ (.A(_06784_),
    .B(_06795_),
    .C(_06938_),
    .Y(_06959_));
 sky130_fd_sc_hd__o21ba_2 _20309_ (.A1(_05777_),
    .A2(_05798_),
    .B1_N(_05766_),
    .X(_06970_));
 sky130_fd_sc_hd__o21ba_2 _20310_ (.A1(_05667_),
    .A2(_05689_),
    .B1_N(_05656_),
    .X(_06981_));
 sky130_fd_sc_hd__and4_2 _20311_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[16]),
    .D(iX[17]),
    .X(_06992_));
 sky130_fd_sc_hd__a22oi_2 _20312_ (.A1(iY[7]),
    .A2(iX[16]),
    .B1(iX[17]),
    .B2(iY[6]),
    .Y(_07003_));
 sky130_fd_sc_hd__nor2_2 _20313_ (.A(_06992_),
    .B(_07003_),
    .Y(_07014_));
 sky130_fd_sc_hd__nand2_2 _20314_ (.A(iY[8]),
    .B(iX[15]),
    .Y(_07025_));
 sky130_fd_sc_hd__xnor2_2 _20315_ (.A(_07014_),
    .B(_07025_),
    .Y(_07036_));
 sky130_fd_sc_hd__xnor2_2 _20316_ (.A(_06981_),
    .B(_07036_),
    .Y(_07047_));
 sky130_fd_sc_hd__xnor2_2 _20317_ (.A(_06970_),
    .B(_07047_),
    .Y(_07058_));
 sky130_fd_sc_hd__nand3_2 _20318_ (.A(_06948_),
    .B(_06959_),
    .C(_07058_),
    .Y(_07069_));
 sky130_fd_sc_hd__a21o_2 _20319_ (.A1(_06948_),
    .A2(_06959_),
    .B1(_07058_),
    .X(_07080_));
 sky130_fd_sc_hd__nand2_2 _20320_ (.A(_05722_),
    .B(_05842_),
    .Y(_07091_));
 sky130_fd_sc_hd__and3_2 _20321_ (.A(_07069_),
    .B(_07080_),
    .C(_07091_),
    .X(_07102_));
 sky130_fd_sc_hd__a21oi_2 _20322_ (.A1(_07069_),
    .A2(_07080_),
    .B1(_07091_),
    .Y(_07113_));
 sky130_fd_sc_hd__and2b_2 _20323_ (.A_N(_06040_),
    .B(_06029_),
    .X(_07124_));
 sky130_fd_sc_hd__or2b_2 _20324_ (.A(_05755_),
    .B_N(_05809_),
    .X(_07135_));
 sky130_fd_sc_hd__or2b_2 _20325_ (.A(_05744_),
    .B_N(_05820_),
    .X(_07146_));
 sky130_fd_sc_hd__and4_2 _20326_ (.A(iX[10]),
    .B(iX[11]),
    .C(iY[12]),
    .D(iY[13]),
    .X(_07157_));
 sky130_fd_sc_hd__a22oi_2 _20327_ (.A1(iX[11]),
    .A2(iY[12]),
    .B1(iY[13]),
    .B2(iX[10]),
    .Y(_07168_));
 sky130_fd_sc_hd__nor2_2 _20328_ (.A(_07157_),
    .B(_07168_),
    .Y(_07179_));
 sky130_fd_sc_hd__nand2_2 _20329_ (.A(iX[9]),
    .B(iY[14]),
    .Y(_07190_));
 sky130_fd_sc_hd__xnor2_2 _20330_ (.A(_07179_),
    .B(_07190_),
    .Y(_07201_));
 sky130_fd_sc_hd__and4_2 _20331_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[13]),
    .D(iX[14]),
    .X(_07211_));
 sky130_fd_sc_hd__a22oi_2 _20332_ (.A1(iY[10]),
    .A2(iX[13]),
    .B1(iX[14]),
    .B2(iY[9]),
    .Y(_07222_));
 sky130_fd_sc_hd__and4bb_2 _20333_ (.A_N(_07211_),
    .B_N(_07222_),
    .C(iY[11]),
    .D(iX[12]),
    .X(_07233_));
 sky130_fd_sc_hd__o2bb2a_2 _20334_ (.A1_N(iY[11]),
    .A2_N(iX[12]),
    .B1(_07211_),
    .B2(_07222_),
    .X(_07244_));
 sky130_fd_sc_hd__nor2_2 _20335_ (.A(_07233_),
    .B(_07244_),
    .Y(_07255_));
 sky130_fd_sc_hd__o21ba_2 _20336_ (.A1(_05996_),
    .A2(_06018_),
    .B1_N(_05985_),
    .X(_07266_));
 sky130_fd_sc_hd__xnor2_2 _20337_ (.A(_07255_),
    .B(_07266_),
    .Y(_07277_));
 sky130_fd_sc_hd__and2_2 _20338_ (.A(_07201_),
    .B(_07277_),
    .X(_07288_));
 sky130_fd_sc_hd__nor2_2 _20339_ (.A(_07201_),
    .B(_07277_),
    .Y(_07299_));
 sky130_fd_sc_hd__or2_2 _20340_ (.A(_07288_),
    .B(_07299_),
    .X(_07310_));
 sky130_fd_sc_hd__a21o_2 _20341_ (.A1(_07135_),
    .A2(_07146_),
    .B1(_07310_),
    .X(_07321_));
 sky130_fd_sc_hd__nand3_2 _20342_ (.A(_07135_),
    .B(_07146_),
    .C(_07310_),
    .Y(_07332_));
 sky130_fd_sc_hd__o211ai_2 _20343_ (.A1(_07124_),
    .A2(_06062_),
    .B1(_07321_),
    .C1(_07332_),
    .Y(_07343_));
 sky130_fd_sc_hd__a211o_2 _20344_ (.A1(_07321_),
    .A2(_07332_),
    .B1(_07124_),
    .C1(_06062_),
    .X(_07354_));
 sky130_fd_sc_hd__and4bb_2 _20345_ (.A_N(_07102_),
    .B_N(_07113_),
    .C(_07343_),
    .D(_07354_),
    .X(_07365_));
 sky130_fd_sc_hd__a2bb2oi_2 _20346_ (.A1_N(_07102_),
    .A2_N(_07113_),
    .B1(_07343_),
    .B2(_07354_),
    .Y(_07376_));
 sky130_fd_sc_hd__a211o_2 _20347_ (.A1(_06773_),
    .A2(_06149_),
    .B1(_07365_),
    .C1(_07376_),
    .X(_07387_));
 sky130_fd_sc_hd__o211ai_2 _20348_ (.A1(_07365_),
    .A2(_07376_),
    .B1(_06773_),
    .C1(_06149_),
    .Y(_07398_));
 sky130_fd_sc_hd__inv_2 _20349_ (.A(_06456_),
    .Y(_07409_));
 sky130_fd_sc_hd__and4_2 _20350_ (.A(iX[1]),
    .B(iX[2]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_07420_));
 sky130_fd_sc_hd__a22o_2 _20351_ (.A1(iX[2]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[1]),
    .X(_07431_));
 sky130_fd_sc_hd__and2b_2 _20352_ (.A_N(_07420_),
    .B(_07431_),
    .X(_07442_));
 sky130_fd_sc_hd__nand2_2 _20353_ (.A(iX[0]),
    .B(iY[23]),
    .Y(_07452_));
 sky130_fd_sc_hd__xnor2_2 _20354_ (.A(_07442_),
    .B(_07452_),
    .Y(_07463_));
 sky130_fd_sc_hd__and4_2 _20355_ (.A(iX[4]),
    .B(iX[5]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_07474_));
 sky130_fd_sc_hd__a22o_2 _20356_ (.A1(iX[5]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[4]),
    .X(_07485_));
 sky130_fd_sc_hd__and2b_2 _20357_ (.A_N(_07474_),
    .B(_07485_),
    .X(_07496_));
 sky130_fd_sc_hd__nand2_2 _20358_ (.A(iX[3]),
    .B(iY[20]),
    .Y(_07507_));
 sky130_fd_sc_hd__xnor2_2 _20359_ (.A(_07496_),
    .B(_07507_),
    .Y(_07518_));
 sky130_fd_sc_hd__a31o_2 _20360_ (.A1(iX[2]),
    .A2(iY[20]),
    .A3(_06237_),
    .B1(_06226_),
    .X(_07529_));
 sky130_fd_sc_hd__xor2_2 _20361_ (.A(_07518_),
    .B(_07529_),
    .X(_07540_));
 sky130_fd_sc_hd__and2_2 _20362_ (.A(_07463_),
    .B(_07540_),
    .X(_07551_));
 sky130_fd_sc_hd__nor2_2 _20363_ (.A(_07463_),
    .B(_07540_),
    .Y(_07562_));
 sky130_fd_sc_hd__or2_2 _20364_ (.A(_07551_),
    .B(_07562_),
    .X(_07573_));
 sky130_fd_sc_hd__or2b_2 _20365_ (.A(_06347_),
    .B_N(_06401_),
    .X(_07584_));
 sky130_fd_sc_hd__nand2_2 _20366_ (.A(_06336_),
    .B(_06412_),
    .Y(_07595_));
 sky130_fd_sc_hd__a31o_2 _20367_ (.A1(iX[5]),
    .A2(iY[17]),
    .A3(_06379_),
    .B1(_06358_),
    .X(_07606_));
 sky130_fd_sc_hd__o21ba_2 _20368_ (.A1(_05941_),
    .A2(_05963_),
    .B1_N(_05930_),
    .X(_07617_));
 sky130_fd_sc_hd__and4_2 _20369_ (.A(iX[7]),
    .B(iX[8]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_07628_));
 sky130_fd_sc_hd__a22oi_2 _20370_ (.A1(iX[8]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[7]),
    .Y(_07639_));
 sky130_fd_sc_hd__and4bb_2 _20371_ (.A_N(_07628_),
    .B_N(_07639_),
    .C(iX[6]),
    .D(iY[17]),
    .X(_07650_));
 sky130_fd_sc_hd__o2bb2a_2 _20372_ (.A1_N(iX[6]),
    .A2_N(iY[17]),
    .B1(_07628_),
    .B2(_07639_),
    .X(_07661_));
 sky130_fd_sc_hd__nor2_2 _20373_ (.A(_07650_),
    .B(_07661_),
    .Y(_07672_));
 sky130_fd_sc_hd__xnor2_2 _20374_ (.A(_07617_),
    .B(_07672_),
    .Y(_07683_));
 sky130_fd_sc_hd__xnor2_2 _20375_ (.A(_07606_),
    .B(_07683_),
    .Y(_07693_));
 sky130_fd_sc_hd__a21oi_2 _20376_ (.A1(_07584_),
    .A2(_07595_),
    .B1(_07693_),
    .Y(_07704_));
 sky130_fd_sc_hd__and3_2 _20377_ (.A(_07584_),
    .B(_07595_),
    .C(_07693_),
    .X(_07715_));
 sky130_fd_sc_hd__or3_2 _20378_ (.A(_07573_),
    .B(_07704_),
    .C(_07715_),
    .X(_07726_));
 sky130_fd_sc_hd__o21ai_2 _20379_ (.A1(_07704_),
    .A2(_07715_),
    .B1(_07573_),
    .Y(_07737_));
 sky130_fd_sc_hd__nand2_2 _20380_ (.A(_07726_),
    .B(_07737_),
    .Y(_07748_));
 sky130_fd_sc_hd__a21oi_2 _20381_ (.A1(_06094_),
    .A2(_06116_),
    .B1(_07748_),
    .Y(_07759_));
 sky130_fd_sc_hd__and3_2 _20382_ (.A(_06094_),
    .B(_06116_),
    .C(_07748_),
    .X(_07770_));
 sky130_fd_sc_hd__a211oi_2 _20383_ (.A1(_06434_),
    .A2(_07409_),
    .B1(_07759_),
    .C1(_07770_),
    .Y(_07781_));
 sky130_fd_sc_hd__o211a_2 _20384_ (.A1(_07759_),
    .A2(_07770_),
    .B1(_06434_),
    .C1(_07409_),
    .X(_07792_));
 sky130_fd_sc_hd__nor2_2 _20385_ (.A(_07781_),
    .B(_07792_),
    .Y(_07803_));
 sky130_fd_sc_hd__nand3_2 _20386_ (.A(_07387_),
    .B(_07398_),
    .C(_07803_),
    .Y(_07814_));
 sky130_fd_sc_hd__a21o_2 _20387_ (.A1(_07387_),
    .A2(_07398_),
    .B1(_07803_),
    .X(_07825_));
 sky130_fd_sc_hd__o211a_2 _20388_ (.A1(_06160_),
    .A2(_06522_),
    .B1(_07814_),
    .C1(_07825_),
    .X(_07836_));
 sky130_fd_sc_hd__a211oi_2 _20389_ (.A1(_07814_),
    .A2(_07825_),
    .B1(_06160_),
    .C1(_06522_),
    .Y(_07847_));
 sky130_fd_sc_hd__nor2_2 _20390_ (.A(_07836_),
    .B(_07847_),
    .Y(_07858_));
 sky130_fd_sc_hd__o21ai_2 _20391_ (.A1(_06182_),
    .A2(_06500_),
    .B1(_06478_),
    .Y(_07869_));
 sky130_fd_sc_hd__inv_2 _20392_ (.A(_06292_),
    .Y(_07880_));
 sky130_fd_sc_hd__and2b_2 _20393_ (.A_N(_06281_),
    .B(_06270_),
    .X(_07891_));
 sky130_fd_sc_hd__nand2_2 _20394_ (.A(_06204_),
    .B(_07891_),
    .Y(_07902_));
 sky130_fd_sc_hd__or2_2 _20395_ (.A(_06204_),
    .B(_07891_),
    .X(_07913_));
 sky130_fd_sc_hd__a2bb2o_2 _20396_ (.A1_N(_06215_),
    .A2_N(_07880_),
    .B1(_07902_),
    .B2(_07913_),
    .X(_07924_));
 sky130_fd_sc_hd__xor2_2 _20397_ (.A(_07869_),
    .B(_07924_),
    .X(_07935_));
 sky130_fd_sc_hd__xnor2_2 _20398_ (.A(_07858_),
    .B(_07935_),
    .Y(_07946_));
 sky130_fd_sc_hd__a21o_2 _20399_ (.A1(_06544_),
    .A2(_06762_),
    .B1(_07946_),
    .X(_07956_));
 sky130_fd_sc_hd__nand3_2 _20400_ (.A(_06544_),
    .B(_06762_),
    .C(_07946_),
    .Y(_07967_));
 sky130_fd_sc_hd__and3_2 _20401_ (.A(_06588_),
    .B(_07956_),
    .C(_07967_),
    .X(_07978_));
 sky130_fd_sc_hd__a21oi_2 _20402_ (.A1(_07956_),
    .A2(_07967_),
    .B1(_06588_),
    .Y(_07989_));
 sky130_fd_sc_hd__or2_2 _20403_ (.A(_07978_),
    .B(_07989_),
    .X(_08000_));
 sky130_fd_sc_hd__nand2_2 _20404_ (.A(_06643_),
    .B(_06654_),
    .Y(_08011_));
 sky130_fd_sc_hd__o21a_2 _20405_ (.A1(_05350_),
    .A2(_06664_),
    .B1(_08011_),
    .X(_08022_));
 sky130_fd_sc_hd__xor2_2 _20406_ (.A(_08000_),
    .B(_08022_),
    .X(_08033_));
 sky130_fd_sc_hd__xor2_2 _20407_ (.A(_06751_),
    .B(_08033_),
    .X(_08044_));
 sky130_fd_sc_hd__o21ba_2 _20408_ (.A1(_06708_),
    .A2(_06730_),
    .B1_N(_06697_),
    .X(_08055_));
 sky130_fd_sc_hd__xor2_2 _20409_ (.A(_08044_),
    .B(_08055_),
    .X(_08066_));
 sky130_fd_sc_hd__inv_2 _20410_ (.A(_08066_),
    .Y(oO[23]));
 sky130_fd_sc_hd__nor2_2 _20411_ (.A(_05448_),
    .B(_05492_),
    .Y(_08087_));
 sky130_fd_sc_hd__nand2_2 _20412_ (.A(_06719_),
    .B(_08044_),
    .Y(_08098_));
 sky130_fd_sc_hd__o21ai_2 _20413_ (.A1(_06751_),
    .A2(_06697_),
    .B1(_08033_),
    .Y(_08109_));
 sky130_fd_sc_hd__o21a_2 _20414_ (.A1(_08087_),
    .A2(_08098_),
    .B1(_08109_),
    .X(_08120_));
 sky130_fd_sc_hd__inv_2 _20415_ (.A(_04265_),
    .Y(_08131_));
 sky130_fd_sc_hd__a2111o_2 _20416_ (.A1(_03146_),
    .A2(_03157_),
    .B1(_08131_),
    .C1(_05470_),
    .D1(_08098_),
    .X(_08142_));
 sky130_fd_sc_hd__nand2_2 _20417_ (.A(_08120_),
    .B(_08142_),
    .Y(_08153_));
 sky130_fd_sc_hd__nor2_2 _20418_ (.A(_08000_),
    .B(_08022_),
    .Y(_08163_));
 sky130_fd_sc_hd__nand2_2 _20419_ (.A(_07869_),
    .B(_07924_),
    .Y(_08174_));
 sky130_fd_sc_hd__inv_2 _20420_ (.A(_07836_),
    .Y(_08185_));
 sky130_fd_sc_hd__nand2_2 _20421_ (.A(_07858_),
    .B(_07935_),
    .Y(_08196_));
 sky130_fd_sc_hd__or2b_2 _20422_ (.A(_06861_),
    .B_N(_06850_),
    .X(_08207_));
 sky130_fd_sc_hd__nand2_2 _20423_ (.A(_06872_),
    .B(_06927_),
    .Y(_08218_));
 sky130_fd_sc_hd__and4_2 _20424_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[23]),
    .D(iX[24]),
    .X(_08229_));
 sky130_fd_sc_hd__a22oi_2 _20425_ (.A1(iY[1]),
    .A2(iX[23]),
    .B1(iX[24]),
    .B2(iY[0]),
    .Y(_08240_));
 sky130_fd_sc_hd__nor2_2 _20426_ (.A(_08229_),
    .B(_08240_),
    .Y(_08251_));
 sky130_fd_sc_hd__nand2_2 _20427_ (.A(iY[2]),
    .B(iX[22]),
    .Y(_08262_));
 sky130_fd_sc_hd__xnor2_2 _20428_ (.A(_08251_),
    .B(_08262_),
    .Y(_08273_));
 sky130_fd_sc_hd__o21ba_2 _20429_ (.A1(_06817_),
    .A2(_06839_),
    .B1_N(_06806_),
    .X(_08284_));
 sky130_fd_sc_hd__xnor2_2 _20430_ (.A(_08273_),
    .B(_08284_),
    .Y(_08295_));
 sky130_fd_sc_hd__and4_2 _20431_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[20]),
    .D(iX[21]),
    .X(_08306_));
 sky130_fd_sc_hd__a22oi_2 _20432_ (.A1(iY[4]),
    .A2(iX[20]),
    .B1(iX[21]),
    .B2(iY[3]),
    .Y(_08317_));
 sky130_fd_sc_hd__nor2_2 _20433_ (.A(_08306_),
    .B(_08317_),
    .Y(_08328_));
 sky130_fd_sc_hd__nand2_2 _20434_ (.A(iY[5]),
    .B(iX[19]),
    .Y(_08339_));
 sky130_fd_sc_hd__xnor2_2 _20435_ (.A(_08328_),
    .B(_08339_),
    .Y(_08350_));
 sky130_fd_sc_hd__xnor2_2 _20436_ (.A(_08295_),
    .B(_08350_),
    .Y(_08361_));
 sky130_fd_sc_hd__a21o_2 _20437_ (.A1(_08207_),
    .A2(_08218_),
    .B1(_08361_),
    .X(_08371_));
 sky130_fd_sc_hd__nand3_2 _20438_ (.A(_08207_),
    .B(_08218_),
    .C(_08361_),
    .Y(_08382_));
 sky130_fd_sc_hd__o21ba_2 _20439_ (.A1(_07003_),
    .A2(_07025_),
    .B1_N(_06992_),
    .X(_08393_));
 sky130_fd_sc_hd__o21ba_2 _20440_ (.A1(_06894_),
    .A2(_06916_),
    .B1_N(_06883_),
    .X(_08404_));
 sky130_fd_sc_hd__and4_2 _20441_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[17]),
    .D(iX[18]),
    .X(_08415_));
 sky130_fd_sc_hd__a22oi_2 _20442_ (.A1(iY[7]),
    .A2(iX[17]),
    .B1(iX[18]),
    .B2(iY[6]),
    .Y(_08426_));
 sky130_fd_sc_hd__nor2_2 _20443_ (.A(_08415_),
    .B(_08426_),
    .Y(_08437_));
 sky130_fd_sc_hd__nand2_2 _20444_ (.A(iY[8]),
    .B(iX[16]),
    .Y(_08448_));
 sky130_fd_sc_hd__xnor2_2 _20445_ (.A(_08437_),
    .B(_08448_),
    .Y(_08459_));
 sky130_fd_sc_hd__xnor2_2 _20446_ (.A(_08404_),
    .B(_08459_),
    .Y(_08470_));
 sky130_fd_sc_hd__xnor2_2 _20447_ (.A(_08393_),
    .B(_08470_),
    .Y(_08481_));
 sky130_fd_sc_hd__and3_2 _20448_ (.A(_08371_),
    .B(_08382_),
    .C(_08481_),
    .X(_08492_));
 sky130_fd_sc_hd__a21oi_2 _20449_ (.A1(_08371_),
    .A2(_08382_),
    .B1(_08481_),
    .Y(_08503_));
 sky130_fd_sc_hd__nor2_2 _20450_ (.A(_08492_),
    .B(_08503_),
    .Y(_08514_));
 sky130_fd_sc_hd__nand2_2 _20451_ (.A(_06948_),
    .B(_07069_),
    .Y(_08525_));
 sky130_fd_sc_hd__xnor2_2 _20452_ (.A(_08514_),
    .B(_08525_),
    .Y(_08536_));
 sky130_fd_sc_hd__and2b_2 _20453_ (.A_N(_07266_),
    .B(_07255_),
    .X(_08547_));
 sky130_fd_sc_hd__or2b_2 _20454_ (.A(_06981_),
    .B_N(_07036_),
    .X(_08557_));
 sky130_fd_sc_hd__or2b_2 _20455_ (.A(_06970_),
    .B_N(_07047_),
    .X(_08568_));
 sky130_fd_sc_hd__and4_2 _20456_ (.A(iX[11]),
    .B(iX[12]),
    .C(iY[12]),
    .D(iY[13]),
    .X(_08579_));
 sky130_fd_sc_hd__a22oi_2 _20457_ (.A1(iX[12]),
    .A2(iY[12]),
    .B1(iY[13]),
    .B2(iX[11]),
    .Y(_08590_));
 sky130_fd_sc_hd__nor2_2 _20458_ (.A(_08579_),
    .B(_08590_),
    .Y(_08601_));
 sky130_fd_sc_hd__nand2_2 _20459_ (.A(iX[10]),
    .B(iY[14]),
    .Y(_08612_));
 sky130_fd_sc_hd__xnor2_2 _20460_ (.A(_08601_),
    .B(_08612_),
    .Y(_08623_));
 sky130_fd_sc_hd__and4_2 _20461_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[14]),
    .D(iX[15]),
    .X(_08634_));
 sky130_fd_sc_hd__a22oi_2 _20462_ (.A1(iY[10]),
    .A2(iX[14]),
    .B1(iX[15]),
    .B2(iY[9]),
    .Y(_08645_));
 sky130_fd_sc_hd__nor2_2 _20463_ (.A(_08634_),
    .B(_08645_),
    .Y(_08656_));
 sky130_fd_sc_hd__nand2_2 _20464_ (.A(iY[11]),
    .B(iX[13]),
    .Y(_08667_));
 sky130_fd_sc_hd__xnor2_2 _20465_ (.A(_08656_),
    .B(_08667_),
    .Y(_08678_));
 sky130_fd_sc_hd__nor2_2 _20466_ (.A(_07211_),
    .B(_07233_),
    .Y(_08689_));
 sky130_fd_sc_hd__xnor2_2 _20467_ (.A(_08678_),
    .B(_08689_),
    .Y(_08700_));
 sky130_fd_sc_hd__xnor2_2 _20468_ (.A(_08623_),
    .B(_08700_),
    .Y(_08711_));
 sky130_fd_sc_hd__a21oi_2 _20469_ (.A1(_08557_),
    .A2(_08568_),
    .B1(_08711_),
    .Y(_08722_));
 sky130_fd_sc_hd__inv_2 _20470_ (.A(_08722_),
    .Y(_08733_));
 sky130_fd_sc_hd__nand3_2 _20471_ (.A(_08557_),
    .B(_08568_),
    .C(_08711_),
    .Y(_08744_));
 sky130_fd_sc_hd__o211a_2 _20472_ (.A1(_08547_),
    .A2(_07288_),
    .B1(_08733_),
    .C1(_08744_),
    .X(_08755_));
 sky130_fd_sc_hd__a211o_2 _20473_ (.A1(_08733_),
    .A2(_08744_),
    .B1(_08547_),
    .C1(_07288_),
    .X(_08765_));
 sky130_fd_sc_hd__or3b_2 _20474_ (.A(_08536_),
    .B(_08755_),
    .C_N(_08765_),
    .X(_08776_));
 sky130_fd_sc_hd__inv_2 _20475_ (.A(_08755_),
    .Y(_08787_));
 sky130_fd_sc_hd__a21bo_2 _20476_ (.A1(_08787_),
    .A2(_08765_),
    .B1_N(_08536_),
    .X(_08798_));
 sky130_fd_sc_hd__o211a_2 _20477_ (.A1(_07102_),
    .A2(_07365_),
    .B1(_08776_),
    .C1(_08798_),
    .X(_08809_));
 sky130_fd_sc_hd__a211oi_2 _20478_ (.A1(_08776_),
    .A2(_08798_),
    .B1(_07102_),
    .C1(_07365_),
    .Y(_08820_));
 sky130_fd_sc_hd__inv_2 _20479_ (.A(_07704_),
    .Y(_08831_));
 sky130_fd_sc_hd__and4_2 _20480_ (.A(iX[2]),
    .B(iX[3]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_08842_));
 sky130_fd_sc_hd__a22oi_2 _20481_ (.A1(iX[3]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[2]),
    .Y(_08853_));
 sky130_fd_sc_hd__nor2_2 _20482_ (.A(_08842_),
    .B(_08853_),
    .Y(_08864_));
 sky130_fd_sc_hd__nand2_2 _20483_ (.A(iX[1]),
    .B(iY[23]),
    .Y(_08875_));
 sky130_fd_sc_hd__xnor2_2 _20484_ (.A(_08864_),
    .B(_08875_),
    .Y(_08886_));
 sky130_fd_sc_hd__and4_2 _20485_ (.A(iX[5]),
    .B(iX[6]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_08897_));
 sky130_fd_sc_hd__a22oi_2 _20486_ (.A1(iX[6]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[5]),
    .Y(_08908_));
 sky130_fd_sc_hd__nor2_2 _20487_ (.A(_08897_),
    .B(_08908_),
    .Y(_08919_));
 sky130_fd_sc_hd__nand2_2 _20488_ (.A(iX[4]),
    .B(iY[20]),
    .Y(_08929_));
 sky130_fd_sc_hd__xnor2_2 _20489_ (.A(_08919_),
    .B(_08929_),
    .Y(_08940_));
 sky130_fd_sc_hd__a31o_2 _20490_ (.A1(iX[3]),
    .A2(iY[20]),
    .A3(_07485_),
    .B1(_07474_),
    .X(_08951_));
 sky130_fd_sc_hd__xor2_2 _20491_ (.A(_08940_),
    .B(_08951_),
    .X(_08962_));
 sky130_fd_sc_hd__and2_2 _20492_ (.A(_08886_),
    .B(_08962_),
    .X(_08973_));
 sky130_fd_sc_hd__nor2_2 _20493_ (.A(_08886_),
    .B(_08962_),
    .Y(_08984_));
 sky130_fd_sc_hd__or2_2 _20494_ (.A(_08973_),
    .B(_08984_),
    .X(_08995_));
 sky130_fd_sc_hd__or3_2 _20495_ (.A(_07617_),
    .B(_07650_),
    .C(_07661_),
    .X(_09006_));
 sky130_fd_sc_hd__nand2_2 _20496_ (.A(_07606_),
    .B(_07683_),
    .Y(_09017_));
 sky130_fd_sc_hd__o21ba_2 _20497_ (.A1(_07168_),
    .A2(_07190_),
    .B1_N(_07157_),
    .X(_09028_));
 sky130_fd_sc_hd__and4_2 _20498_ (.A(iX[8]),
    .B(iX[9]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_09039_));
 sky130_fd_sc_hd__a22oi_2 _20499_ (.A1(iX[9]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[8]),
    .Y(_09050_));
 sky130_fd_sc_hd__and4bb_2 _20500_ (.A_N(_09039_),
    .B_N(_09050_),
    .C(iX[7]),
    .D(iY[17]),
    .X(_09061_));
 sky130_fd_sc_hd__o2bb2a_2 _20501_ (.A1_N(iX[7]),
    .A2_N(iY[17]),
    .B1(_09039_),
    .B2(_09050_),
    .X(_09072_));
 sky130_fd_sc_hd__nor2_2 _20502_ (.A(_09061_),
    .B(_09072_),
    .Y(_09083_));
 sky130_fd_sc_hd__xnor2_2 _20503_ (.A(_09028_),
    .B(_09083_),
    .Y(_09093_));
 sky130_fd_sc_hd__o21ai_2 _20504_ (.A1(_07628_),
    .A2(_07650_),
    .B1(_09093_),
    .Y(_09104_));
 sky130_fd_sc_hd__or3_2 _20505_ (.A(_07628_),
    .B(_07650_),
    .C(_09093_),
    .X(_09115_));
 sky130_fd_sc_hd__nand2_2 _20506_ (.A(_09104_),
    .B(_09115_),
    .Y(_09126_));
 sky130_fd_sc_hd__a21oi_2 _20507_ (.A1(_09006_),
    .A2(_09017_),
    .B1(_09126_),
    .Y(_09137_));
 sky130_fd_sc_hd__and3_2 _20508_ (.A(_09006_),
    .B(_09017_),
    .C(_09126_),
    .X(_09148_));
 sky130_fd_sc_hd__nor3_2 _20509_ (.A(_08995_),
    .B(_09137_),
    .C(_09148_),
    .Y(_09159_));
 sky130_fd_sc_hd__o21a_2 _20510_ (.A1(_09137_),
    .A2(_09148_),
    .B1(_08995_),
    .X(_09170_));
 sky130_fd_sc_hd__a211oi_2 _20511_ (.A1(_07321_),
    .A2(_07343_),
    .B1(_09159_),
    .C1(_09170_),
    .Y(_09181_));
 sky130_fd_sc_hd__o211a_2 _20512_ (.A1(_09159_),
    .A2(_09170_),
    .B1(_07321_),
    .C1(_07343_),
    .X(_09192_));
 sky130_fd_sc_hd__a211oi_2 _20513_ (.A1(_08831_),
    .A2(_07726_),
    .B1(_09181_),
    .C1(_09192_),
    .Y(_09203_));
 sky130_fd_sc_hd__o211a_2 _20514_ (.A1(_09181_),
    .A2(_09192_),
    .B1(_08831_),
    .C1(_07726_),
    .X(_09214_));
 sky130_fd_sc_hd__nor4_2 _20515_ (.A(_08809_),
    .B(_08820_),
    .C(_09203_),
    .D(_09214_),
    .Y(_09225_));
 sky130_fd_sc_hd__o22a_2 _20516_ (.A1(_08809_),
    .A2(_08820_),
    .B1(_09203_),
    .B2(_09214_),
    .X(_09235_));
 sky130_fd_sc_hd__a211oi_2 _20517_ (.A1(_07387_),
    .A2(_07814_),
    .B1(_09225_),
    .C1(_09235_),
    .Y(_09246_));
 sky130_fd_sc_hd__o211a_2 _20518_ (.A1(_09225_),
    .A2(_09235_),
    .B1(_07387_),
    .C1(_07814_),
    .X(_09257_));
 sky130_fd_sc_hd__or2_2 _20519_ (.A(_09246_),
    .B(_09257_),
    .X(_09268_));
 sky130_fd_sc_hd__and2_2 _20520_ (.A(_07518_),
    .B(_07529_),
    .X(_09279_));
 sky130_fd_sc_hd__a31o_2 _20521_ (.A1(iX[0]),
    .A2(iY[23]),
    .A3(_07431_),
    .B1(_07420_),
    .X(_09290_));
 sky130_fd_sc_hd__and3_2 _20522_ (.A(iX[0]),
    .B(iY[24]),
    .C(_09290_),
    .X(_09301_));
 sky130_fd_sc_hd__a21oi_2 _20523_ (.A1(iX[0]),
    .A2(iY[24]),
    .B1(_09290_),
    .Y(_09312_));
 sky130_fd_sc_hd__nor2_2 _20524_ (.A(_09301_),
    .B(_09312_),
    .Y(_09323_));
 sky130_fd_sc_hd__o21ai_2 _20525_ (.A1(_09279_),
    .A2(_07551_),
    .B1(_09323_),
    .Y(_09334_));
 sky130_fd_sc_hd__or3_2 _20526_ (.A(_09279_),
    .B(_07551_),
    .C(_09323_),
    .X(_09345_));
 sky130_fd_sc_hd__and2_2 _20527_ (.A(_09334_),
    .B(_09345_),
    .X(_09356_));
 sky130_fd_sc_hd__xnor2_2 _20528_ (.A(_07902_),
    .B(_09356_),
    .Y(_09367_));
 sky130_fd_sc_hd__o21a_2 _20529_ (.A1(_07759_),
    .A2(_07781_),
    .B1(_09367_),
    .X(_09378_));
 sky130_fd_sc_hd__nor3_2 _20530_ (.A(_07759_),
    .B(_07781_),
    .C(_09367_),
    .Y(_09389_));
 sky130_fd_sc_hd__or2_2 _20531_ (.A(_09378_),
    .B(_09389_),
    .X(_09399_));
 sky130_fd_sc_hd__xnor2_2 _20532_ (.A(_09268_),
    .B(_09399_),
    .Y(_09410_));
 sky130_fd_sc_hd__a21oi_2 _20533_ (.A1(_08185_),
    .A2(_08196_),
    .B1(_09410_),
    .Y(_09421_));
 sky130_fd_sc_hd__and3_2 _20534_ (.A(_08185_),
    .B(_08196_),
    .C(_09410_),
    .X(_09432_));
 sky130_fd_sc_hd__nor3_2 _20535_ (.A(_08174_),
    .B(_09421_),
    .C(_09432_),
    .Y(_09443_));
 sky130_fd_sc_hd__o21a_2 _20536_ (.A1(_09421_),
    .A2(_09432_),
    .B1(_08174_),
    .X(_09454_));
 sky130_fd_sc_hd__nor2_2 _20537_ (.A(_09443_),
    .B(_09454_),
    .Y(_09465_));
 sky130_fd_sc_hd__a21bo_2 _20538_ (.A1(_06588_),
    .A2(_07967_),
    .B1_N(_07956_),
    .X(_09476_));
 sky130_fd_sc_hd__xor2_2 _20539_ (.A(_09465_),
    .B(_09476_),
    .X(_09487_));
 sky130_fd_sc_hd__and2_2 _20540_ (.A(_08163_),
    .B(_09487_),
    .X(_09498_));
 sky130_fd_sc_hd__nor2_2 _20541_ (.A(_08163_),
    .B(_09487_),
    .Y(_09509_));
 sky130_fd_sc_hd__nor2_2 _20542_ (.A(_09498_),
    .B(_09509_),
    .Y(_09520_));
 sky130_fd_sc_hd__xnor2_2 _20543_ (.A(_08153_),
    .B(_09520_),
    .Y(_09530_));
 sky130_fd_sc_hd__inv_2 _20544_ (.A(_09530_),
    .Y(oO[24]));
 sky130_fd_sc_hd__and2_2 _20545_ (.A(_09465_),
    .B(_09476_),
    .X(_09551_));
 sky130_fd_sc_hd__nor2_2 _20546_ (.A(_09268_),
    .B(_09399_),
    .Y(_09562_));
 sky130_fd_sc_hd__a21oi_2 _20547_ (.A1(_08207_),
    .A2(_08218_),
    .B1(_08361_),
    .Y(_09573_));
 sky130_fd_sc_hd__or2b_2 _20548_ (.A(_08284_),
    .B_N(_08273_),
    .X(_09584_));
 sky130_fd_sc_hd__nand2_2 _20549_ (.A(_08295_),
    .B(_08350_),
    .Y(_09595_));
 sky130_fd_sc_hd__and4_2 _20550_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[24]),
    .D(iX[25]),
    .X(_09606_));
 sky130_fd_sc_hd__a22oi_2 _20551_ (.A1(iY[1]),
    .A2(iX[24]),
    .B1(iX[25]),
    .B2(iY[0]),
    .Y(_09617_));
 sky130_fd_sc_hd__nor2_2 _20552_ (.A(_09606_),
    .B(_09617_),
    .Y(_09628_));
 sky130_fd_sc_hd__nand2_2 _20553_ (.A(iY[2]),
    .B(iX[23]),
    .Y(_09639_));
 sky130_fd_sc_hd__xnor2_2 _20554_ (.A(_09628_),
    .B(_09639_),
    .Y(_09649_));
 sky130_fd_sc_hd__o21ba_2 _20555_ (.A1(_08240_),
    .A2(_08262_),
    .B1_N(_08229_),
    .X(_09660_));
 sky130_fd_sc_hd__xnor2_2 _20556_ (.A(_09649_),
    .B(_09660_),
    .Y(_09671_));
 sky130_fd_sc_hd__and4_2 _20557_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[21]),
    .D(iX[22]),
    .X(_09682_));
 sky130_fd_sc_hd__a22oi_2 _20558_ (.A1(iY[4]),
    .A2(iX[21]),
    .B1(iX[22]),
    .B2(iY[3]),
    .Y(_09693_));
 sky130_fd_sc_hd__nor2_2 _20559_ (.A(_09682_),
    .B(_09693_),
    .Y(_09704_));
 sky130_fd_sc_hd__nand2_2 _20560_ (.A(iY[5]),
    .B(iX[20]),
    .Y(_09715_));
 sky130_fd_sc_hd__xnor2_2 _20561_ (.A(_09704_),
    .B(_09715_),
    .Y(_09725_));
 sky130_fd_sc_hd__nand2_2 _20562_ (.A(_09671_),
    .B(_09725_),
    .Y(_09736_));
 sky130_fd_sc_hd__or2_2 _20563_ (.A(_09671_),
    .B(_09725_),
    .X(_09747_));
 sky130_fd_sc_hd__nand2_2 _20564_ (.A(_09736_),
    .B(_09747_),
    .Y(_09758_));
 sky130_fd_sc_hd__a21o_2 _20565_ (.A1(_09584_),
    .A2(_09595_),
    .B1(_09758_),
    .X(_09769_));
 sky130_fd_sc_hd__nand3_2 _20566_ (.A(_09584_),
    .B(_09595_),
    .C(_09758_),
    .Y(_09780_));
 sky130_fd_sc_hd__o21ba_2 _20567_ (.A1(_08426_),
    .A2(_08448_),
    .B1_N(_08415_),
    .X(_09791_));
 sky130_fd_sc_hd__o21ba_2 _20568_ (.A1(_08317_),
    .A2(_08339_),
    .B1_N(_08306_),
    .X(_09801_));
 sky130_fd_sc_hd__and4_2 _20569_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[18]),
    .D(iX[19]),
    .X(_09812_));
 sky130_fd_sc_hd__a22oi_2 _20570_ (.A1(iY[7]),
    .A2(iX[18]),
    .B1(iX[19]),
    .B2(iY[6]),
    .Y(_09823_));
 sky130_fd_sc_hd__nor2_2 _20571_ (.A(_09812_),
    .B(_09823_),
    .Y(_09834_));
 sky130_fd_sc_hd__nand2_2 _20572_ (.A(iY[8]),
    .B(iX[17]),
    .Y(_09845_));
 sky130_fd_sc_hd__xnor2_2 _20573_ (.A(_09834_),
    .B(_09845_),
    .Y(_09856_));
 sky130_fd_sc_hd__xnor2_2 _20574_ (.A(_09801_),
    .B(_09856_),
    .Y(_09867_));
 sky130_fd_sc_hd__xnor2_2 _20575_ (.A(_09791_),
    .B(_09867_),
    .Y(_09877_));
 sky130_fd_sc_hd__nand3_2 _20576_ (.A(_09769_),
    .B(_09780_),
    .C(_09877_),
    .Y(_09888_));
 sky130_fd_sc_hd__a21o_2 _20577_ (.A1(_09769_),
    .A2(_09780_),
    .B1(_09877_),
    .X(_09899_));
 sky130_fd_sc_hd__o211a_2 _20578_ (.A1(_09573_),
    .A2(_08492_),
    .B1(_09888_),
    .C1(_09899_),
    .X(_09910_));
 sky130_fd_sc_hd__a211oi_2 _20579_ (.A1(_09888_),
    .A2(_09899_),
    .B1(_09573_),
    .C1(_08492_),
    .Y(_09921_));
 sky130_fd_sc_hd__or2_2 _20580_ (.A(_09910_),
    .B(_09921_),
    .X(_09931_));
 sky130_fd_sc_hd__and2b_2 _20581_ (.A_N(_08689_),
    .B(_08678_),
    .X(_09942_));
 sky130_fd_sc_hd__a21o_2 _20582_ (.A1(_08623_),
    .A2(_08700_),
    .B1(_09942_),
    .X(_09953_));
 sky130_fd_sc_hd__or2b_2 _20583_ (.A(_08404_),
    .B_N(_08459_),
    .X(_09963_));
 sky130_fd_sc_hd__or2b_2 _20584_ (.A(_08393_),
    .B_N(_08470_),
    .X(_09974_));
 sky130_fd_sc_hd__and4_2 _20585_ (.A(iX[12]),
    .B(iY[12]),
    .C(iX[13]),
    .D(iY[13]),
    .X(_09985_));
 sky130_fd_sc_hd__a22oi_2 _20586_ (.A1(iY[12]),
    .A2(iX[13]),
    .B1(iY[13]),
    .B2(iX[12]),
    .Y(_09996_));
 sky130_fd_sc_hd__nor2_2 _20587_ (.A(_09985_),
    .B(_09996_),
    .Y(_10006_));
 sky130_fd_sc_hd__nand2_2 _20588_ (.A(iX[11]),
    .B(iY[14]),
    .Y(_10016_));
 sky130_fd_sc_hd__xnor2_2 _20589_ (.A(_10006_),
    .B(_10016_),
    .Y(_10025_));
 sky130_fd_sc_hd__and4_2 _20590_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[15]),
    .D(iX[16]),
    .X(_10035_));
 sky130_fd_sc_hd__a22oi_2 _20591_ (.A1(iY[10]),
    .A2(iX[15]),
    .B1(iX[16]),
    .B2(iY[9]),
    .Y(_10043_));
 sky130_fd_sc_hd__and4bb_2 _20592_ (.A_N(_10035_),
    .B_N(_10043_),
    .C(iY[11]),
    .D(iX[14]),
    .X(_10053_));
 sky130_fd_sc_hd__o2bb2a_2 _20593_ (.A1_N(iY[11]),
    .A2_N(iX[14]),
    .B1(_10035_),
    .B2(_10043_),
    .X(_10062_));
 sky130_fd_sc_hd__nor2_2 _20594_ (.A(_10053_),
    .B(_10062_),
    .Y(_10072_));
 sky130_fd_sc_hd__o21ba_2 _20595_ (.A1(_08645_),
    .A2(_08667_),
    .B1_N(_08634_),
    .X(_10081_));
 sky130_fd_sc_hd__xnor2_2 _20596_ (.A(_10072_),
    .B(_10081_),
    .Y(_10090_));
 sky130_fd_sc_hd__and2_2 _20597_ (.A(_10025_),
    .B(_10090_),
    .X(_10100_));
 sky130_fd_sc_hd__nor2_2 _20598_ (.A(_10025_),
    .B(_10090_),
    .Y(_10108_));
 sky130_fd_sc_hd__or2_2 _20599_ (.A(_10100_),
    .B(_10108_),
    .X(_10118_));
 sky130_fd_sc_hd__a21o_2 _20600_ (.A1(_09963_),
    .A2(_09974_),
    .B1(_10118_),
    .X(_10127_));
 sky130_fd_sc_hd__nand3_2 _20601_ (.A(_09963_),
    .B(_09974_),
    .C(_10118_),
    .Y(_10137_));
 sky130_fd_sc_hd__nand3_2 _20602_ (.A(_09953_),
    .B(_10127_),
    .C(_10137_),
    .Y(_10145_));
 sky130_fd_sc_hd__a21o_2 _20603_ (.A1(_10127_),
    .A2(_10137_),
    .B1(_09953_),
    .X(_10155_));
 sky130_fd_sc_hd__nand2_2 _20604_ (.A(_10145_),
    .B(_10155_),
    .Y(_10163_));
 sky130_fd_sc_hd__xor2_2 _20605_ (.A(_09931_),
    .B(_10163_),
    .X(_10167_));
 sky130_fd_sc_hd__a21bo_2 _20606_ (.A1(_08514_),
    .A2(_08525_),
    .B1_N(_08776_),
    .X(_10168_));
 sky130_fd_sc_hd__xnor2_2 _20607_ (.A(_10167_),
    .B(_10168_),
    .Y(_10169_));
 sky130_fd_sc_hd__and4_2 _20608_ (.A(iX[3]),
    .B(iX[4]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_10170_));
 sky130_fd_sc_hd__a22oi_2 _20609_ (.A1(iX[4]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[3]),
    .Y(_10171_));
 sky130_fd_sc_hd__nor2_2 _20610_ (.A(_10170_),
    .B(_10171_),
    .Y(_10172_));
 sky130_fd_sc_hd__nand2_2 _20611_ (.A(iX[2]),
    .B(iY[23]),
    .Y(_10173_));
 sky130_fd_sc_hd__xnor2_2 _20612_ (.A(_10172_),
    .B(_10173_),
    .Y(_10174_));
 sky130_fd_sc_hd__and4_2 _20613_ (.A(iX[6]),
    .B(iX[7]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_10175_));
 sky130_fd_sc_hd__a22oi_2 _20614_ (.A1(iX[7]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[6]),
    .Y(_10176_));
 sky130_fd_sc_hd__nor2_2 _20615_ (.A(_10175_),
    .B(_10176_),
    .Y(_10177_));
 sky130_fd_sc_hd__nand2_2 _20616_ (.A(iX[5]),
    .B(iY[20]),
    .Y(_10178_));
 sky130_fd_sc_hd__xnor2_2 _20617_ (.A(_10177_),
    .B(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__o21ba_2 _20618_ (.A1(_08908_),
    .A2(_08929_),
    .B1_N(_08897_),
    .X(_10180_));
 sky130_fd_sc_hd__xnor2_2 _20619_ (.A(_10179_),
    .B(_10180_),
    .Y(_10181_));
 sky130_fd_sc_hd__nand2_2 _20620_ (.A(_10174_),
    .B(_10181_),
    .Y(_10182_));
 sky130_fd_sc_hd__or2_2 _20621_ (.A(_10174_),
    .B(_10181_),
    .X(_10183_));
 sky130_fd_sc_hd__nand2_2 _20622_ (.A(_10182_),
    .B(_10183_),
    .Y(_10184_));
 sky130_fd_sc_hd__or3_2 _20623_ (.A(_09028_),
    .B(_09061_),
    .C(_09072_),
    .X(_10185_));
 sky130_fd_sc_hd__o21ba_2 _20624_ (.A1(_08590_),
    .A2(_08612_),
    .B1_N(_08579_),
    .X(_10186_));
 sky130_fd_sc_hd__and4_2 _20625_ (.A(iX[9]),
    .B(iX[10]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_10187_));
 sky130_fd_sc_hd__a22oi_2 _20626_ (.A1(iX[10]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[9]),
    .Y(_10188_));
 sky130_fd_sc_hd__and4bb_2 _20627_ (.A_N(_10187_),
    .B_N(_10188_),
    .C(iX[8]),
    .D(iY[17]),
    .X(_10189_));
 sky130_fd_sc_hd__o2bb2a_2 _20628_ (.A1_N(iX[8]),
    .A2_N(iY[17]),
    .B1(_10187_),
    .B2(_10188_),
    .X(_10190_));
 sky130_fd_sc_hd__nor2_2 _20629_ (.A(_10189_),
    .B(_10190_),
    .Y(_10191_));
 sky130_fd_sc_hd__xnor2_2 _20630_ (.A(_10186_),
    .B(_10191_),
    .Y(_10192_));
 sky130_fd_sc_hd__o21ai_2 _20631_ (.A1(_09039_),
    .A2(_09061_),
    .B1(_10192_),
    .Y(_10193_));
 sky130_fd_sc_hd__or3_2 _20632_ (.A(_09039_),
    .B(_09061_),
    .C(_10192_),
    .X(_10194_));
 sky130_fd_sc_hd__nand2_2 _20633_ (.A(_10193_),
    .B(_10194_),
    .Y(_10195_));
 sky130_fd_sc_hd__a21oi_2 _20634_ (.A1(_10185_),
    .A2(_09104_),
    .B1(_10195_),
    .Y(_10196_));
 sky130_fd_sc_hd__and3_2 _20635_ (.A(_10185_),
    .B(_09104_),
    .C(_10195_),
    .X(_10197_));
 sky130_fd_sc_hd__or3_2 _20636_ (.A(_10184_),
    .B(_10196_),
    .C(_10197_),
    .X(_10198_));
 sky130_fd_sc_hd__o21ai_2 _20637_ (.A1(_10196_),
    .A2(_10197_),
    .B1(_10184_),
    .Y(_10199_));
 sky130_fd_sc_hd__o211a_2 _20638_ (.A1(_08722_),
    .A2(_08755_),
    .B1(_10198_),
    .C1(_10199_),
    .X(_10200_));
 sky130_fd_sc_hd__inv_2 _20639_ (.A(_10200_),
    .Y(_10201_));
 sky130_fd_sc_hd__a211o_2 _20640_ (.A1(_10198_),
    .A2(_10199_),
    .B1(_08722_),
    .C1(_08755_),
    .X(_10202_));
 sky130_fd_sc_hd__o211a_2 _20641_ (.A1(_09137_),
    .A2(_09159_),
    .B1(_10201_),
    .C1(_10202_),
    .X(_10203_));
 sky130_fd_sc_hd__a211oi_2 _20642_ (.A1(_10201_),
    .A2(_10202_),
    .B1(_09137_),
    .C1(_09159_),
    .Y(_10204_));
 sky130_fd_sc_hd__nor2_2 _20643_ (.A(_10203_),
    .B(_10204_),
    .Y(_10205_));
 sky130_fd_sc_hd__xnor2_2 _20644_ (.A(_10169_),
    .B(_10205_),
    .Y(_10206_));
 sky130_fd_sc_hd__o21a_2 _20645_ (.A1(_08809_),
    .A2(_09225_),
    .B1(_10206_),
    .X(_10207_));
 sky130_fd_sc_hd__nor3_2 _20646_ (.A(_08809_),
    .B(_09225_),
    .C(_10206_),
    .Y(_10208_));
 sky130_fd_sc_hd__and3_2 _20647_ (.A(_06204_),
    .B(_07891_),
    .C(_09356_),
    .X(_10209_));
 sky130_fd_sc_hd__and2_2 _20648_ (.A(_08940_),
    .B(_08951_),
    .X(_10210_));
 sky130_fd_sc_hd__a31o_2 _20649_ (.A1(iX[1]),
    .A2(iY[23]),
    .A3(_08864_),
    .B1(_08842_),
    .X(_10211_));
 sky130_fd_sc_hd__a22o_2 _20650_ (.A1(iX[1]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[0]),
    .X(_10212_));
 sky130_fd_sc_hd__and4_2 _20651_ (.A(iX[0]),
    .B(iX[1]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_10213_));
 sky130_fd_sc_hd__inv_2 _20652_ (.A(_10213_),
    .Y(_10214_));
 sky130_fd_sc_hd__and3_2 _20653_ (.A(_10211_),
    .B(_10212_),
    .C(_10214_),
    .X(_10215_));
 sky130_fd_sc_hd__a21oi_2 _20654_ (.A1(_10212_),
    .A2(_10214_),
    .B1(_10211_),
    .Y(_10216_));
 sky130_fd_sc_hd__nor2_2 _20655_ (.A(_10215_),
    .B(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__o21ai_2 _20656_ (.A1(_10210_),
    .A2(_08973_),
    .B1(_10217_),
    .Y(_10218_));
 sky130_fd_sc_hd__or3_2 _20657_ (.A(_10210_),
    .B(_08973_),
    .C(_10217_),
    .X(_10219_));
 sky130_fd_sc_hd__and2_2 _20658_ (.A(_10218_),
    .B(_10219_),
    .X(_10220_));
 sky130_fd_sc_hd__nand2_2 _20659_ (.A(_09301_),
    .B(_10220_),
    .Y(_10221_));
 sky130_fd_sc_hd__or2_2 _20660_ (.A(_09301_),
    .B(_10220_),
    .X(_10222_));
 sky130_fd_sc_hd__nand2_2 _20661_ (.A(_10221_),
    .B(_10222_),
    .Y(_10223_));
 sky130_fd_sc_hd__nor2_2 _20662_ (.A(_09334_),
    .B(_10223_),
    .Y(_10224_));
 sky130_fd_sc_hd__and2_2 _20663_ (.A(_09334_),
    .B(_10223_),
    .X(_10225_));
 sky130_fd_sc_hd__nor2_2 _20664_ (.A(_10224_),
    .B(_10225_),
    .Y(_10226_));
 sky130_fd_sc_hd__o21a_2 _20665_ (.A1(_09181_),
    .A2(_09203_),
    .B1(_10226_),
    .X(_10227_));
 sky130_fd_sc_hd__nor3_2 _20666_ (.A(_09181_),
    .B(_09203_),
    .C(_10226_),
    .Y(_10228_));
 sky130_fd_sc_hd__nor2_2 _20667_ (.A(_10227_),
    .B(_10228_),
    .Y(_10229_));
 sky130_fd_sc_hd__xnor2_2 _20668_ (.A(_10209_),
    .B(_10229_),
    .Y(_10230_));
 sky130_fd_sc_hd__nor3_2 _20669_ (.A(_10207_),
    .B(_10208_),
    .C(_10230_),
    .Y(_10231_));
 sky130_fd_sc_hd__o21a_2 _20670_ (.A1(_10207_),
    .A2(_10208_),
    .B1(_10230_),
    .X(_10232_));
 sky130_fd_sc_hd__nor2_2 _20671_ (.A(_10231_),
    .B(_10232_),
    .Y(_10233_));
 sky130_fd_sc_hd__o21ai_2 _20672_ (.A1(_09246_),
    .A2(_09562_),
    .B1(_10233_),
    .Y(_10234_));
 sky130_fd_sc_hd__or3_2 _20673_ (.A(_09246_),
    .B(_09562_),
    .C(_10233_),
    .X(_10235_));
 sky130_fd_sc_hd__nand3_2 _20674_ (.A(_09378_),
    .B(_10234_),
    .C(_10235_),
    .Y(_10236_));
 sky130_fd_sc_hd__a21o_2 _20675_ (.A1(_10234_),
    .A2(_10235_),
    .B1(_09378_),
    .X(_10237_));
 sky130_fd_sc_hd__o211ai_2 _20676_ (.A1(_09421_),
    .A2(_09443_),
    .B1(_10236_),
    .C1(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__a211o_2 _20677_ (.A1(_10236_),
    .A2(_10237_),
    .B1(_09421_),
    .C1(_09443_),
    .X(_10239_));
 sky130_fd_sc_hd__and3_2 _20678_ (.A(_09551_),
    .B(_10238_),
    .C(_10239_),
    .X(_10240_));
 sky130_fd_sc_hd__a21oi_2 _20679_ (.A1(_10238_),
    .A2(_10239_),
    .B1(_09551_),
    .Y(_10241_));
 sky130_fd_sc_hd__nor2_2 _20680_ (.A(_10240_),
    .B(_10241_),
    .Y(_10242_));
 sky130_fd_sc_hd__a21oi_2 _20681_ (.A1(_08153_),
    .A2(_09520_),
    .B1(_09498_),
    .Y(_10243_));
 sky130_fd_sc_hd__xnor2_2 _20682_ (.A(_10242_),
    .B(_10243_),
    .Y(oO[25]));
 sky130_fd_sc_hd__nand2_2 _20683_ (.A(_09520_),
    .B(_10242_),
    .Y(_10244_));
 sky130_fd_sc_hd__a21o_2 _20684_ (.A1(_08120_),
    .A2(_08142_),
    .B1(_10244_),
    .X(_10245_));
 sky130_fd_sc_hd__a21oi_2 _20685_ (.A1(_09498_),
    .A2(_10242_),
    .B1(_10240_),
    .Y(_10246_));
 sky130_fd_sc_hd__nand2_2 _20686_ (.A(_10167_),
    .B(_10168_),
    .Y(_10247_));
 sky130_fd_sc_hd__or3_2 _20687_ (.A(_10169_),
    .B(_10203_),
    .C(_10204_),
    .X(_10248_));
 sky130_fd_sc_hd__nor2_2 _20688_ (.A(_09931_),
    .B(_10163_),
    .Y(_10249_));
 sky130_fd_sc_hd__or2b_2 _20689_ (.A(_09660_),
    .B_N(_09649_),
    .X(_10250_));
 sky130_fd_sc_hd__and4_2 _20690_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[25]),
    .D(iX[26]),
    .X(_10251_));
 sky130_fd_sc_hd__a22oi_2 _20691_ (.A1(iY[1]),
    .A2(iX[25]),
    .B1(iX[26]),
    .B2(iY[0]),
    .Y(_10252_));
 sky130_fd_sc_hd__nor2_2 _20692_ (.A(_10251_),
    .B(_10252_),
    .Y(_10253_));
 sky130_fd_sc_hd__nand2_2 _20693_ (.A(iY[2]),
    .B(iX[24]),
    .Y(_10254_));
 sky130_fd_sc_hd__xnor2_2 _20694_ (.A(_10253_),
    .B(_10254_),
    .Y(_10255_));
 sky130_fd_sc_hd__o21ba_2 _20695_ (.A1(_09617_),
    .A2(_09639_),
    .B1_N(_09606_),
    .X(_10256_));
 sky130_fd_sc_hd__xnor2_2 _20696_ (.A(_10255_),
    .B(_10256_),
    .Y(_10257_));
 sky130_fd_sc_hd__and4_2 _20697_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[22]),
    .D(iX[23]),
    .X(_10258_));
 sky130_fd_sc_hd__a22oi_2 _20698_ (.A1(iY[4]),
    .A2(iX[22]),
    .B1(iX[23]),
    .B2(iY[3]),
    .Y(_10259_));
 sky130_fd_sc_hd__nor2_2 _20699_ (.A(_10258_),
    .B(_10259_),
    .Y(_10260_));
 sky130_fd_sc_hd__nand2_2 _20700_ (.A(iY[5]),
    .B(iX[21]),
    .Y(_10261_));
 sky130_fd_sc_hd__xnor2_2 _20701_ (.A(_10260_),
    .B(_10261_),
    .Y(_10262_));
 sky130_fd_sc_hd__nand2_2 _20702_ (.A(_10257_),
    .B(_10262_),
    .Y(_10263_));
 sky130_fd_sc_hd__or2_2 _20703_ (.A(_10257_),
    .B(_10262_),
    .X(_10264_));
 sky130_fd_sc_hd__nand2_2 _20704_ (.A(_10263_),
    .B(_10264_),
    .Y(_10265_));
 sky130_fd_sc_hd__a21o_2 _20705_ (.A1(_10250_),
    .A2(_09736_),
    .B1(_10265_),
    .X(_10266_));
 sky130_fd_sc_hd__nand3_2 _20706_ (.A(_10250_),
    .B(_09736_),
    .C(_10265_),
    .Y(_10267_));
 sky130_fd_sc_hd__o21ba_2 _20707_ (.A1(_09823_),
    .A2(_09845_),
    .B1_N(_09812_),
    .X(_10268_));
 sky130_fd_sc_hd__o21ba_2 _20708_ (.A1(_09693_),
    .A2(_09715_),
    .B1_N(_09682_),
    .X(_10269_));
 sky130_fd_sc_hd__and4_2 _20709_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[19]),
    .D(iX[20]),
    .X(_10270_));
 sky130_fd_sc_hd__a22oi_2 _20710_ (.A1(iY[7]),
    .A2(iX[19]),
    .B1(iX[20]),
    .B2(iY[6]),
    .Y(_10271_));
 sky130_fd_sc_hd__nor2_2 _20711_ (.A(_10270_),
    .B(_10271_),
    .Y(_10272_));
 sky130_fd_sc_hd__nand2_2 _20712_ (.A(iY[8]),
    .B(iX[18]),
    .Y(_10273_));
 sky130_fd_sc_hd__xnor2_2 _20713_ (.A(_10272_),
    .B(_10273_),
    .Y(_10274_));
 sky130_fd_sc_hd__xnor2_2 _20714_ (.A(_10269_),
    .B(_10274_),
    .Y(_10275_));
 sky130_fd_sc_hd__xnor2_2 _20715_ (.A(_10268_),
    .B(_10275_),
    .Y(_10276_));
 sky130_fd_sc_hd__and3_2 _20716_ (.A(_10266_),
    .B(_10267_),
    .C(_10276_),
    .X(_10277_));
 sky130_fd_sc_hd__a21oi_2 _20717_ (.A1(_10266_),
    .A2(_10267_),
    .B1(_10276_),
    .Y(_10278_));
 sky130_fd_sc_hd__nor2_2 _20718_ (.A(_10277_),
    .B(_10278_),
    .Y(_10279_));
 sky130_fd_sc_hd__nand2_2 _20719_ (.A(_09769_),
    .B(_09888_),
    .Y(_10280_));
 sky130_fd_sc_hd__xnor2_2 _20720_ (.A(_10279_),
    .B(_10280_),
    .Y(_10281_));
 sky130_fd_sc_hd__and2b_2 _20721_ (.A_N(_10081_),
    .B(_10072_),
    .X(_10282_));
 sky130_fd_sc_hd__or2b_2 _20722_ (.A(_09801_),
    .B_N(_09856_),
    .X(_10283_));
 sky130_fd_sc_hd__or2b_2 _20723_ (.A(_09791_),
    .B_N(_09867_),
    .X(_10284_));
 sky130_fd_sc_hd__and4_2 _20724_ (.A(iY[12]),
    .B(iX[13]),
    .C(iY[13]),
    .D(iX[14]),
    .X(_10285_));
 sky130_fd_sc_hd__a22oi_2 _20725_ (.A1(iX[13]),
    .A2(iY[13]),
    .B1(iX[14]),
    .B2(iY[12]),
    .Y(_10286_));
 sky130_fd_sc_hd__nor2_2 _20726_ (.A(_10285_),
    .B(_10286_),
    .Y(_10287_));
 sky130_fd_sc_hd__nand2_2 _20727_ (.A(iX[12]),
    .B(iY[14]),
    .Y(_10288_));
 sky130_fd_sc_hd__xnor2_2 _20728_ (.A(_10287_),
    .B(_10288_),
    .Y(_10289_));
 sky130_fd_sc_hd__and4_2 _20729_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[16]),
    .D(iX[17]),
    .X(_10290_));
 sky130_fd_sc_hd__a22oi_2 _20730_ (.A1(iY[10]),
    .A2(iX[16]),
    .B1(iX[17]),
    .B2(iY[9]),
    .Y(_10291_));
 sky130_fd_sc_hd__nor2_2 _20731_ (.A(_10290_),
    .B(_10291_),
    .Y(_10292_));
 sky130_fd_sc_hd__nand2_2 _20732_ (.A(iY[11]),
    .B(iX[15]),
    .Y(_10293_));
 sky130_fd_sc_hd__xnor2_2 _20733_ (.A(_10292_),
    .B(_10293_),
    .Y(_10294_));
 sky130_fd_sc_hd__o21ai_2 _20734_ (.A1(_10035_),
    .A2(_10053_),
    .B1(_10294_),
    .Y(_10295_));
 sky130_fd_sc_hd__or3_2 _20735_ (.A(_10035_),
    .B(_10053_),
    .C(_10294_),
    .X(_10296_));
 sky130_fd_sc_hd__and2_2 _20736_ (.A(_10295_),
    .B(_10296_),
    .X(_10297_));
 sky130_fd_sc_hd__xnor2_2 _20737_ (.A(_10289_),
    .B(_10297_),
    .Y(_10298_));
 sky130_fd_sc_hd__a21oi_2 _20738_ (.A1(_10283_),
    .A2(_10284_),
    .B1(_10298_),
    .Y(_10299_));
 sky130_fd_sc_hd__inv_2 _20739_ (.A(_10299_),
    .Y(_10300_));
 sky130_fd_sc_hd__nand3_2 _20740_ (.A(_10283_),
    .B(_10284_),
    .C(_10298_),
    .Y(_10301_));
 sky130_fd_sc_hd__o211a_2 _20741_ (.A1(_10282_),
    .A2(_10100_),
    .B1(_10300_),
    .C1(_10301_),
    .X(_10302_));
 sky130_fd_sc_hd__a211o_2 _20742_ (.A1(_10300_),
    .A2(_10301_),
    .B1(_10282_),
    .C1(_10100_),
    .X(_10303_));
 sky130_fd_sc_hd__or3b_2 _20743_ (.A(_10281_),
    .B(_10302_),
    .C_N(_10303_),
    .X(_10304_));
 sky130_fd_sc_hd__inv_2 _20744_ (.A(_10302_),
    .Y(_10305_));
 sky130_fd_sc_hd__a21bo_2 _20745_ (.A1(_10305_),
    .A2(_10303_),
    .B1_N(_10281_),
    .X(_10306_));
 sky130_fd_sc_hd__o211a_2 _20746_ (.A1(_09910_),
    .A2(_10249_),
    .B1(_10304_),
    .C1(_10306_),
    .X(_10307_));
 sky130_fd_sc_hd__a211oi_2 _20747_ (.A1(_10304_),
    .A2(_10306_),
    .B1(_09910_),
    .C1(_10249_),
    .Y(_10308_));
 sky130_fd_sc_hd__a21o_2 _20748_ (.A1(_10185_),
    .A2(_09104_),
    .B1(_10195_),
    .X(_10309_));
 sky130_fd_sc_hd__and4_2 _20749_ (.A(iX[4]),
    .B(iX[5]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_10310_));
 sky130_fd_sc_hd__a22oi_2 _20750_ (.A1(iX[5]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[4]),
    .Y(_10311_));
 sky130_fd_sc_hd__nor2_2 _20751_ (.A(_10310_),
    .B(_10311_),
    .Y(_10312_));
 sky130_fd_sc_hd__nand2_2 _20752_ (.A(iX[3]),
    .B(iY[23]),
    .Y(_10313_));
 sky130_fd_sc_hd__xnor2_2 _20753_ (.A(_10312_),
    .B(_10313_),
    .Y(_10314_));
 sky130_fd_sc_hd__and4_2 _20754_ (.A(iX[7]),
    .B(iX[8]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_10315_));
 sky130_fd_sc_hd__a22oi_2 _20755_ (.A1(iX[8]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[7]),
    .Y(_10316_));
 sky130_fd_sc_hd__nor2_2 _20756_ (.A(_10315_),
    .B(_10316_),
    .Y(_10317_));
 sky130_fd_sc_hd__nand2_2 _20757_ (.A(iX[6]),
    .B(iY[20]),
    .Y(_10318_));
 sky130_fd_sc_hd__xnor2_2 _20758_ (.A(_10317_),
    .B(_10318_),
    .Y(_10319_));
 sky130_fd_sc_hd__o21ba_2 _20759_ (.A1(_10176_),
    .A2(_10178_),
    .B1_N(_10175_),
    .X(_10320_));
 sky130_fd_sc_hd__xnor2_2 _20760_ (.A(_10319_),
    .B(_10320_),
    .Y(_10321_));
 sky130_fd_sc_hd__and2_2 _20761_ (.A(_10314_),
    .B(_10321_),
    .X(_10322_));
 sky130_fd_sc_hd__nor2_2 _20762_ (.A(_10314_),
    .B(_10321_),
    .Y(_10323_));
 sky130_fd_sc_hd__or2_2 _20763_ (.A(_10322_),
    .B(_10323_),
    .X(_10324_));
 sky130_fd_sc_hd__or3_2 _20764_ (.A(_10186_),
    .B(_10189_),
    .C(_10190_),
    .X(_10325_));
 sky130_fd_sc_hd__o21ba_2 _20765_ (.A1(_09996_),
    .A2(_10016_),
    .B1_N(_09985_),
    .X(_10326_));
 sky130_fd_sc_hd__and4_2 _20766_ (.A(iX[10]),
    .B(iX[11]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_10327_));
 sky130_fd_sc_hd__a22oi_2 _20767_ (.A1(iX[11]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[10]),
    .Y(_10328_));
 sky130_fd_sc_hd__and4bb_2 _20768_ (.A_N(_10327_),
    .B_N(_10328_),
    .C(iX[9]),
    .D(iY[17]),
    .X(_10329_));
 sky130_fd_sc_hd__o2bb2a_2 _20769_ (.A1_N(iX[9]),
    .A2_N(iY[17]),
    .B1(_10327_),
    .B2(_10328_),
    .X(_10330_));
 sky130_fd_sc_hd__nor2_2 _20770_ (.A(_10329_),
    .B(_10330_),
    .Y(_10331_));
 sky130_fd_sc_hd__xnor2_2 _20771_ (.A(_10326_),
    .B(_10331_),
    .Y(_10332_));
 sky130_fd_sc_hd__o21ai_2 _20772_ (.A1(_10187_),
    .A2(_10189_),
    .B1(_10332_),
    .Y(_10333_));
 sky130_fd_sc_hd__or3_2 _20773_ (.A(_10187_),
    .B(_10189_),
    .C(_10332_),
    .X(_10334_));
 sky130_fd_sc_hd__nand2_2 _20774_ (.A(_10333_),
    .B(_10334_),
    .Y(_10335_));
 sky130_fd_sc_hd__a21oi_2 _20775_ (.A1(_10325_),
    .A2(_10193_),
    .B1(_10335_),
    .Y(_10336_));
 sky130_fd_sc_hd__and3_2 _20776_ (.A(_10325_),
    .B(_10193_),
    .C(_10335_),
    .X(_10337_));
 sky130_fd_sc_hd__nor3_2 _20777_ (.A(_10324_),
    .B(_10336_),
    .C(_10337_),
    .Y(_10338_));
 sky130_fd_sc_hd__o21a_2 _20778_ (.A1(_10336_),
    .A2(_10337_),
    .B1(_10324_),
    .X(_10339_));
 sky130_fd_sc_hd__a211oi_2 _20779_ (.A1(_10127_),
    .A2(_10145_),
    .B1(_10338_),
    .C1(_10339_),
    .Y(_10340_));
 sky130_fd_sc_hd__o211a_2 _20780_ (.A1(_10338_),
    .A2(_10339_),
    .B1(_10127_),
    .C1(_10145_),
    .X(_10341_));
 sky130_fd_sc_hd__a211oi_2 _20781_ (.A1(_10309_),
    .A2(_10198_),
    .B1(_10340_),
    .C1(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__o211a_2 _20782_ (.A1(_10340_),
    .A2(_10341_),
    .B1(_10309_),
    .C1(_10198_),
    .X(_10343_));
 sky130_fd_sc_hd__nor4_2 _20783_ (.A(_10307_),
    .B(_10308_),
    .C(_10342_),
    .D(_10343_),
    .Y(_10344_));
 sky130_fd_sc_hd__o22a_2 _20784_ (.A1(_10307_),
    .A2(_10308_),
    .B1(_10342_),
    .B2(_10343_),
    .X(_10345_));
 sky130_fd_sc_hd__a211oi_2 _20785_ (.A1(_10247_),
    .A2(_10248_),
    .B1(_10344_),
    .C1(_10345_),
    .Y(_10346_));
 sky130_fd_sc_hd__o211a_2 _20786_ (.A1(_10344_),
    .A2(_10345_),
    .B1(_10247_),
    .C1(_10248_),
    .X(_10347_));
 sky130_fd_sc_hd__or2_2 _20787_ (.A(_10200_),
    .B(_10203_),
    .X(_10348_));
 sky130_fd_sc_hd__or2b_2 _20788_ (.A(_10180_),
    .B_N(_10179_),
    .X(_10349_));
 sky130_fd_sc_hd__o21ba_2 _20789_ (.A1(_10171_),
    .A2(_10173_),
    .B1_N(_10170_),
    .X(_10350_));
 sky130_fd_sc_hd__and4_2 _20790_ (.A(iX[1]),
    .B(iX[2]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_10351_));
 sky130_fd_sc_hd__a22oi_2 _20791_ (.A1(iX[2]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[1]),
    .Y(_10352_));
 sky130_fd_sc_hd__nor2_2 _20792_ (.A(_10351_),
    .B(_10352_),
    .Y(_10353_));
 sky130_fd_sc_hd__nand2_2 _20793_ (.A(iX[0]),
    .B(iY[26]),
    .Y(_10354_));
 sky130_fd_sc_hd__xnor2_2 _20794_ (.A(_10353_),
    .B(_10354_),
    .Y(_10355_));
 sky130_fd_sc_hd__xnor2_2 _20795_ (.A(_10350_),
    .B(_10355_),
    .Y(_10356_));
 sky130_fd_sc_hd__xnor2_2 _20796_ (.A(_10213_),
    .B(_10356_),
    .Y(_10357_));
 sky130_fd_sc_hd__a21oi_2 _20797_ (.A1(_10349_),
    .A2(_10182_),
    .B1(_10357_),
    .Y(_10358_));
 sky130_fd_sc_hd__and3_2 _20798_ (.A(_10349_),
    .B(_10182_),
    .C(_10357_),
    .X(_10359_));
 sky130_fd_sc_hd__nor2_2 _20799_ (.A(_10358_),
    .B(_10359_),
    .Y(_10360_));
 sky130_fd_sc_hd__xnor2_2 _20800_ (.A(_10215_),
    .B(_10360_),
    .Y(_10361_));
 sky130_fd_sc_hd__a21o_2 _20801_ (.A1(_10218_),
    .A2(_10221_),
    .B1(_10361_),
    .X(_10362_));
 sky130_fd_sc_hd__nand3_2 _20802_ (.A(_10218_),
    .B(_10221_),
    .C(_10361_),
    .Y(_10363_));
 sky130_fd_sc_hd__nand2_2 _20803_ (.A(_10362_),
    .B(_10363_),
    .Y(_10364_));
 sky130_fd_sc_hd__xnor2_2 _20804_ (.A(_10348_),
    .B(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__nor2_2 _20805_ (.A(_10224_),
    .B(_10365_),
    .Y(_10366_));
 sky130_fd_sc_hd__and2_2 _20806_ (.A(_10224_),
    .B(_10365_),
    .X(_10367_));
 sky130_fd_sc_hd__or2_2 _20807_ (.A(_10366_),
    .B(_10367_),
    .X(_10368_));
 sky130_fd_sc_hd__or3_2 _20808_ (.A(_10346_),
    .B(_10347_),
    .C(_10368_),
    .X(_10369_));
 sky130_fd_sc_hd__o21ai_2 _20809_ (.A1(_10346_),
    .A2(_10347_),
    .B1(_10368_),
    .Y(_10370_));
 sky130_fd_sc_hd__o211ai_2 _20810_ (.A1(_10207_),
    .A2(_10231_),
    .B1(_10369_),
    .C1(_10370_),
    .Y(_10371_));
 sky130_fd_sc_hd__a211o_2 _20811_ (.A1(_10369_),
    .A2(_10370_),
    .B1(_10207_),
    .C1(_10231_),
    .X(_10372_));
 sky130_fd_sc_hd__nand2_2 _20812_ (.A(_10371_),
    .B(_10372_),
    .Y(_10373_));
 sky130_fd_sc_hd__a21oi_2 _20813_ (.A1(_10209_),
    .A2(_10229_),
    .B1(_10227_),
    .Y(_10374_));
 sky130_fd_sc_hd__xnor2_2 _20814_ (.A(_10373_),
    .B(_10374_),
    .Y(_10375_));
 sky130_fd_sc_hd__a21oi_2 _20815_ (.A1(_10234_),
    .A2(_10236_),
    .B1(_10375_),
    .Y(_10376_));
 sky130_fd_sc_hd__and3_2 _20816_ (.A(_10234_),
    .B(_10236_),
    .C(_10375_),
    .X(_10377_));
 sky130_fd_sc_hd__nor2_2 _20817_ (.A(_10376_),
    .B(_10377_),
    .Y(_10378_));
 sky130_fd_sc_hd__xor2_2 _20818_ (.A(_10238_),
    .B(_10378_),
    .X(_10379_));
 sky130_fd_sc_hd__a21oi_2 _20819_ (.A1(_10245_),
    .A2(_10246_),
    .B1(_10379_),
    .Y(_10380_));
 sky130_fd_sc_hd__and3_2 _20820_ (.A(_10245_),
    .B(_10379_),
    .C(_10246_),
    .X(_10381_));
 sky130_fd_sc_hd__or2_2 _20821_ (.A(_10380_),
    .B(_10381_),
    .X(_10382_));
 sky130_fd_sc_hd__inv_2 _20822_ (.A(_10382_),
    .Y(oO[26]));
 sky130_fd_sc_hd__inv_2 _20823_ (.A(_10371_),
    .Y(_10383_));
 sky130_fd_sc_hd__nor2_2 _20824_ (.A(_10373_),
    .B(_10374_),
    .Y(_10384_));
 sky130_fd_sc_hd__and3_2 _20825_ (.A(_10348_),
    .B(_10362_),
    .C(_10363_),
    .X(_10385_));
 sky130_fd_sc_hd__inv_2 _20826_ (.A(_10369_),
    .Y(_10386_));
 sky130_fd_sc_hd__or2b_2 _20827_ (.A(_10256_),
    .B_N(_10255_),
    .X(_10387_));
 sky130_fd_sc_hd__and4_2 _20828_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[26]),
    .D(iX[27]),
    .X(_10388_));
 sky130_fd_sc_hd__a22oi_2 _20829_ (.A1(iY[1]),
    .A2(iX[26]),
    .B1(iX[27]),
    .B2(iY[0]),
    .Y(_10389_));
 sky130_fd_sc_hd__nor2_2 _20830_ (.A(_10388_),
    .B(_10389_),
    .Y(_10390_));
 sky130_fd_sc_hd__nand2_2 _20831_ (.A(iY[2]),
    .B(iX[25]),
    .Y(_10391_));
 sky130_fd_sc_hd__xnor2_2 _20832_ (.A(_10390_),
    .B(_10391_),
    .Y(_10392_));
 sky130_fd_sc_hd__o21ba_2 _20833_ (.A1(_10252_),
    .A2(_10254_),
    .B1_N(_10251_),
    .X(_10393_));
 sky130_fd_sc_hd__xnor2_2 _20834_ (.A(_10392_),
    .B(_10393_),
    .Y(_10394_));
 sky130_fd_sc_hd__and4_2 _20835_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[23]),
    .D(iX[24]),
    .X(_10395_));
 sky130_fd_sc_hd__a22oi_2 _20836_ (.A1(iY[4]),
    .A2(iX[23]),
    .B1(iX[24]),
    .B2(iY[3]),
    .Y(_10396_));
 sky130_fd_sc_hd__nor2_2 _20837_ (.A(_10395_),
    .B(_10396_),
    .Y(_10397_));
 sky130_fd_sc_hd__nand2_2 _20838_ (.A(iY[5]),
    .B(iX[22]),
    .Y(_10398_));
 sky130_fd_sc_hd__xnor2_2 _20839_ (.A(_10397_),
    .B(_10398_),
    .Y(_10399_));
 sky130_fd_sc_hd__xnor2_2 _20840_ (.A(_10394_),
    .B(_10399_),
    .Y(_10400_));
 sky130_fd_sc_hd__a21o_2 _20841_ (.A1(_10387_),
    .A2(_10263_),
    .B1(_10400_),
    .X(_10401_));
 sky130_fd_sc_hd__nand3_2 _20842_ (.A(_10387_),
    .B(_10263_),
    .C(_10400_),
    .Y(_10402_));
 sky130_fd_sc_hd__o21ba_2 _20843_ (.A1(_10271_),
    .A2(_10273_),
    .B1_N(_10270_),
    .X(_10403_));
 sky130_fd_sc_hd__o21ba_2 _20844_ (.A1(_10259_),
    .A2(_10261_),
    .B1_N(_10258_),
    .X(_10404_));
 sky130_fd_sc_hd__and4_2 _20845_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[20]),
    .D(iX[21]),
    .X(_10405_));
 sky130_fd_sc_hd__a22oi_2 _20846_ (.A1(iY[7]),
    .A2(iX[20]),
    .B1(iX[21]),
    .B2(iY[6]),
    .Y(_10406_));
 sky130_fd_sc_hd__nor2_2 _20847_ (.A(_10405_),
    .B(_10406_),
    .Y(_10407_));
 sky130_fd_sc_hd__nand2_2 _20848_ (.A(iY[8]),
    .B(iX[19]),
    .Y(_10408_));
 sky130_fd_sc_hd__xnor2_2 _20849_ (.A(_10407_),
    .B(_10408_),
    .Y(_10409_));
 sky130_fd_sc_hd__xnor2_2 _20850_ (.A(_10404_),
    .B(_10409_),
    .Y(_10410_));
 sky130_fd_sc_hd__xnor2_2 _20851_ (.A(_10403_),
    .B(_10410_),
    .Y(_10411_));
 sky130_fd_sc_hd__nand3_2 _20852_ (.A(_10401_),
    .B(_10402_),
    .C(_10411_),
    .Y(_10412_));
 sky130_fd_sc_hd__a21o_2 _20853_ (.A1(_10401_),
    .A2(_10402_),
    .B1(_10411_),
    .X(_10413_));
 sky130_fd_sc_hd__nand2_2 _20854_ (.A(_10412_),
    .B(_10413_),
    .Y(_10414_));
 sky130_fd_sc_hd__a21bo_2 _20855_ (.A1(_10267_),
    .A2(_10276_),
    .B1_N(_10266_),
    .X(_10415_));
 sky130_fd_sc_hd__xor2_2 _20856_ (.A(_10414_),
    .B(_10415_),
    .X(_10416_));
 sky130_fd_sc_hd__a21bo_2 _20857_ (.A1(_10289_),
    .A2(_10297_),
    .B1_N(_10295_),
    .X(_10417_));
 sky130_fd_sc_hd__or2b_2 _20858_ (.A(_10269_),
    .B_N(_10274_),
    .X(_10418_));
 sky130_fd_sc_hd__or2b_2 _20859_ (.A(_10268_),
    .B_N(_10275_),
    .X(_10419_));
 sky130_fd_sc_hd__and4_2 _20860_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[14]),
    .D(iX[15]),
    .X(_10420_));
 sky130_fd_sc_hd__a22oi_2 _20861_ (.A1(iY[13]),
    .A2(iX[14]),
    .B1(iX[15]),
    .B2(iY[12]),
    .Y(_10421_));
 sky130_fd_sc_hd__nor2_2 _20862_ (.A(_10420_),
    .B(_10421_),
    .Y(_10422_));
 sky130_fd_sc_hd__nand2_2 _20863_ (.A(iX[13]),
    .B(iY[14]),
    .Y(_10423_));
 sky130_fd_sc_hd__xnor2_2 _20864_ (.A(_10422_),
    .B(_10423_),
    .Y(_10424_));
 sky130_fd_sc_hd__and4_2 _20865_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[17]),
    .D(iX[18]),
    .X(_10425_));
 sky130_fd_sc_hd__a22oi_2 _20866_ (.A1(iY[10]),
    .A2(iX[17]),
    .B1(iX[18]),
    .B2(iY[9]),
    .Y(_10426_));
 sky130_fd_sc_hd__nor2_2 _20867_ (.A(_10425_),
    .B(_10426_),
    .Y(_10427_));
 sky130_fd_sc_hd__nand2_2 _20868_ (.A(iY[11]),
    .B(iX[16]),
    .Y(_10428_));
 sky130_fd_sc_hd__xnor2_2 _20869_ (.A(_10427_),
    .B(_10428_),
    .Y(_10429_));
 sky130_fd_sc_hd__o21ba_2 _20870_ (.A1(_10291_),
    .A2(_10293_),
    .B1_N(_10290_),
    .X(_10430_));
 sky130_fd_sc_hd__xnor2_2 _20871_ (.A(_10429_),
    .B(_10430_),
    .Y(_10431_));
 sky130_fd_sc_hd__and2_2 _20872_ (.A(_10424_),
    .B(_10431_),
    .X(_10432_));
 sky130_fd_sc_hd__nor2_2 _20873_ (.A(_10424_),
    .B(_10431_),
    .Y(_10433_));
 sky130_fd_sc_hd__or2_2 _20874_ (.A(_10432_),
    .B(_10433_),
    .X(_10434_));
 sky130_fd_sc_hd__a21o_2 _20875_ (.A1(_10418_),
    .A2(_10419_),
    .B1(_10434_),
    .X(_10435_));
 sky130_fd_sc_hd__and3_2 _20876_ (.A(_10418_),
    .B(_10419_),
    .C(_10434_),
    .X(_10436_));
 sky130_fd_sc_hd__inv_2 _20877_ (.A(_10436_),
    .Y(_10437_));
 sky130_fd_sc_hd__nand3_2 _20878_ (.A(_10417_),
    .B(_10435_),
    .C(_10437_),
    .Y(_10438_));
 sky130_fd_sc_hd__a21o_2 _20879_ (.A1(_10435_),
    .A2(_10437_),
    .B1(_10417_),
    .X(_10439_));
 sky130_fd_sc_hd__nand2_2 _20880_ (.A(_10438_),
    .B(_10439_),
    .Y(_10440_));
 sky130_fd_sc_hd__nor2_2 _20881_ (.A(_10416_),
    .B(_10440_),
    .Y(_10441_));
 sky130_fd_sc_hd__and2_2 _20882_ (.A(_10416_),
    .B(_10440_),
    .X(_10442_));
 sky130_fd_sc_hd__nor2_2 _20883_ (.A(_10441_),
    .B(_10442_),
    .Y(_10443_));
 sky130_fd_sc_hd__a21bo_2 _20884_ (.A1(_10279_),
    .A2(_10280_),
    .B1_N(_10304_),
    .X(_10444_));
 sky130_fd_sc_hd__xnor2_2 _20885_ (.A(_10443_),
    .B(_10444_),
    .Y(_10445_));
 sky130_fd_sc_hd__and4_2 _20886_ (.A(iX[5]),
    .B(iX[6]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_10446_));
 sky130_fd_sc_hd__a22oi_2 _20887_ (.A1(iX[6]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[5]),
    .Y(_10447_));
 sky130_fd_sc_hd__nor2_2 _20888_ (.A(_10446_),
    .B(_10447_),
    .Y(_10448_));
 sky130_fd_sc_hd__nand2_2 _20889_ (.A(iX[4]),
    .B(iY[23]),
    .Y(_10449_));
 sky130_fd_sc_hd__xnor2_2 _20890_ (.A(_10448_),
    .B(_10449_),
    .Y(_10450_));
 sky130_fd_sc_hd__and4_2 _20891_ (.A(iX[8]),
    .B(iX[9]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_10451_));
 sky130_fd_sc_hd__a22oi_2 _20892_ (.A1(iX[9]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[8]),
    .Y(_10452_));
 sky130_fd_sc_hd__nor2_2 _20893_ (.A(_10451_),
    .B(_10452_),
    .Y(_10453_));
 sky130_fd_sc_hd__nand2_2 _20894_ (.A(iX[7]),
    .B(iY[20]),
    .Y(_10454_));
 sky130_fd_sc_hd__xnor2_2 _20895_ (.A(_10453_),
    .B(_10454_),
    .Y(_10455_));
 sky130_fd_sc_hd__o21ba_2 _20896_ (.A1(_10316_),
    .A2(_10318_),
    .B1_N(_10315_),
    .X(_10456_));
 sky130_fd_sc_hd__xnor2_2 _20897_ (.A(_10455_),
    .B(_10456_),
    .Y(_10457_));
 sky130_fd_sc_hd__and2_2 _20898_ (.A(_10450_),
    .B(_10457_),
    .X(_10458_));
 sky130_fd_sc_hd__nor2_2 _20899_ (.A(_10450_),
    .B(_10457_),
    .Y(_10459_));
 sky130_fd_sc_hd__or2_2 _20900_ (.A(_10458_),
    .B(_10459_),
    .X(_10460_));
 sky130_fd_sc_hd__or3_2 _20901_ (.A(_10326_),
    .B(_10329_),
    .C(_10330_),
    .X(_10461_));
 sky130_fd_sc_hd__o21ba_2 _20902_ (.A1(_10286_),
    .A2(_10288_),
    .B1_N(_10285_),
    .X(_10462_));
 sky130_fd_sc_hd__and4_2 _20903_ (.A(iX[11]),
    .B(iX[12]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_10463_));
 sky130_fd_sc_hd__a22oi_2 _20904_ (.A1(iX[12]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[11]),
    .Y(_10464_));
 sky130_fd_sc_hd__and4bb_2 _20905_ (.A_N(_10463_),
    .B_N(_10464_),
    .C(iX[10]),
    .D(iY[17]),
    .X(_10465_));
 sky130_fd_sc_hd__o2bb2a_2 _20906_ (.A1_N(iX[10]),
    .A2_N(iY[17]),
    .B1(_10463_),
    .B2(_10464_),
    .X(_10466_));
 sky130_fd_sc_hd__nor2_2 _20907_ (.A(_10465_),
    .B(_10466_),
    .Y(_10467_));
 sky130_fd_sc_hd__xnor2_2 _20908_ (.A(_10462_),
    .B(_10467_),
    .Y(_10468_));
 sky130_fd_sc_hd__o21ai_2 _20909_ (.A1(_10327_),
    .A2(_10329_),
    .B1(_10468_),
    .Y(_10469_));
 sky130_fd_sc_hd__or3_2 _20910_ (.A(_10327_),
    .B(_10329_),
    .C(_10468_),
    .X(_10470_));
 sky130_fd_sc_hd__nand2_2 _20911_ (.A(_10469_),
    .B(_10470_),
    .Y(_10471_));
 sky130_fd_sc_hd__a21oi_2 _20912_ (.A1(_10461_),
    .A2(_10333_),
    .B1(_10471_),
    .Y(_10472_));
 sky130_fd_sc_hd__and3_2 _20913_ (.A(_10461_),
    .B(_10333_),
    .C(_10471_),
    .X(_10473_));
 sky130_fd_sc_hd__or3_2 _20914_ (.A(_10460_),
    .B(_10472_),
    .C(_10473_),
    .X(_10474_));
 sky130_fd_sc_hd__o21ai_2 _20915_ (.A1(_10472_),
    .A2(_10473_),
    .B1(_10460_),
    .Y(_10475_));
 sky130_fd_sc_hd__o211a_2 _20916_ (.A1(_10299_),
    .A2(_10302_),
    .B1(_10474_),
    .C1(_10475_),
    .X(_10476_));
 sky130_fd_sc_hd__inv_2 _20917_ (.A(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__a211o_2 _20918_ (.A1(_10474_),
    .A2(_10475_),
    .B1(_10299_),
    .C1(_10302_),
    .X(_10478_));
 sky130_fd_sc_hd__o211a_2 _20919_ (.A1(_10336_),
    .A2(_10338_),
    .B1(_10477_),
    .C1(_10478_),
    .X(_10479_));
 sky130_fd_sc_hd__a211oi_2 _20920_ (.A1(_10477_),
    .A2(_10478_),
    .B1(_10336_),
    .C1(_10338_),
    .Y(_10480_));
 sky130_fd_sc_hd__or3_2 _20921_ (.A(_10445_),
    .B(_10479_),
    .C(_10480_),
    .X(_10481_));
 sky130_fd_sc_hd__o21ai_2 _20922_ (.A1(_10479_),
    .A2(_10480_),
    .B1(_10445_),
    .Y(_10482_));
 sky130_fd_sc_hd__and2_2 _20923_ (.A(_10481_),
    .B(_10482_),
    .X(_10483_));
 sky130_fd_sc_hd__o21ai_2 _20924_ (.A1(_10307_),
    .A2(_10344_),
    .B1(_10483_),
    .Y(_10484_));
 sky130_fd_sc_hd__or3_2 _20925_ (.A(_10307_),
    .B(_10344_),
    .C(_10483_),
    .X(_10485_));
 sky130_fd_sc_hd__and2b_2 _20926_ (.A_N(_10320_),
    .B(_10319_),
    .X(_10486_));
 sky130_fd_sc_hd__o21ba_2 _20927_ (.A1(_10352_),
    .A2(_10354_),
    .B1_N(_10351_),
    .X(_10487_));
 sky130_fd_sc_hd__o21ba_2 _20928_ (.A1(_10311_),
    .A2(_10313_),
    .B1_N(_10310_),
    .X(_10488_));
 sky130_fd_sc_hd__and4_2 _20929_ (.A(iX[2]),
    .B(iX[3]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_10489_));
 sky130_fd_sc_hd__a22oi_2 _20930_ (.A1(iX[3]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[2]),
    .Y(_10490_));
 sky130_fd_sc_hd__nor2_2 _20931_ (.A(_10489_),
    .B(_10490_),
    .Y(_10491_));
 sky130_fd_sc_hd__nand2_2 _20932_ (.A(iX[1]),
    .B(iY[26]),
    .Y(_10492_));
 sky130_fd_sc_hd__xnor2_2 _20933_ (.A(_10491_),
    .B(_10492_),
    .Y(_10493_));
 sky130_fd_sc_hd__xnor2_2 _20934_ (.A(_10488_),
    .B(_10493_),
    .Y(_10494_));
 sky130_fd_sc_hd__xnor2_2 _20935_ (.A(_10487_),
    .B(_10494_),
    .Y(_10495_));
 sky130_fd_sc_hd__o21a_2 _20936_ (.A1(_10486_),
    .A2(_10322_),
    .B1(_10495_),
    .X(_10496_));
 sky130_fd_sc_hd__nor3_2 _20937_ (.A(_10486_),
    .B(_10322_),
    .C(_10495_),
    .Y(_10497_));
 sky130_fd_sc_hd__and2b_2 _20938_ (.A_N(_10350_),
    .B(_10355_),
    .X(_10498_));
 sky130_fd_sc_hd__a21oi_2 _20939_ (.A1(_10213_),
    .A2(_10356_),
    .B1(_10498_),
    .Y(_10499_));
 sky130_fd_sc_hd__nor3_2 _20940_ (.A(_10496_),
    .B(_10497_),
    .C(_10499_),
    .Y(_10500_));
 sky130_fd_sc_hd__o21a_2 _20941_ (.A1(_10496_),
    .A2(_10497_),
    .B1(_10499_),
    .X(_10501_));
 sky130_fd_sc_hd__or2_2 _20942_ (.A(_10500_),
    .B(_10501_),
    .X(_10502_));
 sky130_fd_sc_hd__a21oi_2 _20943_ (.A1(_10215_),
    .A2(_10360_),
    .B1(_10358_),
    .Y(_10503_));
 sky130_fd_sc_hd__or2_2 _20944_ (.A(_10502_),
    .B(_10503_),
    .X(_10504_));
 sky130_fd_sc_hd__nand2_2 _20945_ (.A(_10502_),
    .B(_10503_),
    .Y(_10505_));
 sky130_fd_sc_hd__nand2_2 _20946_ (.A(_10504_),
    .B(_10505_),
    .Y(_10506_));
 sky130_fd_sc_hd__nand2_2 _20947_ (.A(iX[0]),
    .B(iY[27]),
    .Y(_10507_));
 sky130_fd_sc_hd__or2_2 _20948_ (.A(_10506_),
    .B(_10507_),
    .X(_10508_));
 sky130_fd_sc_hd__nand2_2 _20949_ (.A(_10506_),
    .B(_10507_),
    .Y(_10509_));
 sky130_fd_sc_hd__and2_2 _20950_ (.A(_10508_),
    .B(_10509_),
    .X(_10510_));
 sky130_fd_sc_hd__o21a_2 _20951_ (.A1(_10340_),
    .A2(_10342_),
    .B1(_10510_),
    .X(_10511_));
 sky130_fd_sc_hd__nor3_2 _20952_ (.A(_10340_),
    .B(_10342_),
    .C(_10510_),
    .Y(_10512_));
 sky130_fd_sc_hd__o21ai_2 _20953_ (.A1(_10511_),
    .A2(_10512_),
    .B1(_10362_),
    .Y(_10513_));
 sky130_fd_sc_hd__or3_2 _20954_ (.A(_10362_),
    .B(_10511_),
    .C(_10512_),
    .X(_10514_));
 sky130_fd_sc_hd__nand4_2 _20955_ (.A(_10484_),
    .B(_10485_),
    .C(_10513_),
    .D(_10514_),
    .Y(_10515_));
 sky130_fd_sc_hd__a22o_2 _20956_ (.A1(_10484_),
    .A2(_10485_),
    .B1(_10513_),
    .B2(_10514_),
    .X(_10516_));
 sky130_fd_sc_hd__o211ai_2 _20957_ (.A1(_10346_),
    .A2(_10386_),
    .B1(_10515_),
    .C1(_10516_),
    .Y(_10517_));
 sky130_fd_sc_hd__a211o_2 _20958_ (.A1(_10515_),
    .A2(_10516_),
    .B1(_10346_),
    .C1(_10386_),
    .X(_10518_));
 sky130_fd_sc_hd__o211ai_2 _20959_ (.A1(_10385_),
    .A2(_10367_),
    .B1(_10517_),
    .C1(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__a211o_2 _20960_ (.A1(_10517_),
    .A2(_10518_),
    .B1(_10385_),
    .C1(_10367_),
    .X(_10520_));
 sky130_fd_sc_hd__o211ai_2 _20961_ (.A1(_10383_),
    .A2(_10384_),
    .B1(_10519_),
    .C1(_10520_),
    .Y(_10521_));
 sky130_fd_sc_hd__a211o_2 _20962_ (.A1(_10519_),
    .A2(_10520_),
    .B1(_10383_),
    .C1(_10384_),
    .X(_10522_));
 sky130_fd_sc_hd__and3_2 _20963_ (.A(_10376_),
    .B(_10521_),
    .C(_10522_),
    .X(_10523_));
 sky130_fd_sc_hd__a21o_2 _20964_ (.A1(_10521_),
    .A2(_10522_),
    .B1(_10376_),
    .X(_10524_));
 sky130_fd_sc_hd__and2b_2 _20965_ (.A_N(_10523_),
    .B(_10524_),
    .X(_10525_));
 sky130_fd_sc_hd__and2b_2 _20966_ (.A_N(_10238_),
    .B(_10378_),
    .X(_10526_));
 sky130_fd_sc_hd__nor2_2 _20967_ (.A(_10526_),
    .B(_10380_),
    .Y(_10527_));
 sky130_fd_sc_hd__xnor2_2 _20968_ (.A(_10525_),
    .B(_10527_),
    .Y(oO[27]));
 sky130_fd_sc_hd__inv_2 _20969_ (.A(_10511_),
    .Y(_10528_));
 sky130_fd_sc_hd__and3_2 _20970_ (.A(_10412_),
    .B(_10413_),
    .C(_10415_),
    .X(_10529_));
 sky130_fd_sc_hd__or2b_2 _20971_ (.A(_10393_),
    .B_N(_10392_),
    .X(_10530_));
 sky130_fd_sc_hd__nand2_2 _20972_ (.A(_10394_),
    .B(_10399_),
    .Y(_10531_));
 sky130_fd_sc_hd__and4_2 _20973_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[27]),
    .D(iX[28]),
    .X(_10532_));
 sky130_fd_sc_hd__a22oi_2 _20974_ (.A1(iY[1]),
    .A2(iX[27]),
    .B1(iX[28]),
    .B2(iY[0]),
    .Y(_10533_));
 sky130_fd_sc_hd__nor2_2 _20975_ (.A(_10532_),
    .B(_10533_),
    .Y(_10534_));
 sky130_fd_sc_hd__nand2_2 _20976_ (.A(iY[2]),
    .B(iX[26]),
    .Y(_10535_));
 sky130_fd_sc_hd__xnor2_2 _20977_ (.A(_10534_),
    .B(_10535_),
    .Y(_10536_));
 sky130_fd_sc_hd__o21ba_2 _20978_ (.A1(_10389_),
    .A2(_10391_),
    .B1_N(_10388_),
    .X(_10537_));
 sky130_fd_sc_hd__xnor2_2 _20979_ (.A(_10536_),
    .B(_10537_),
    .Y(_10538_));
 sky130_fd_sc_hd__and4_2 _20980_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[24]),
    .D(iX[25]),
    .X(_10539_));
 sky130_fd_sc_hd__a22oi_2 _20981_ (.A1(iY[4]),
    .A2(iX[24]),
    .B1(iX[25]),
    .B2(iY[3]),
    .Y(_10540_));
 sky130_fd_sc_hd__nor2_2 _20982_ (.A(_10539_),
    .B(_10540_),
    .Y(_10541_));
 sky130_fd_sc_hd__nand2_2 _20983_ (.A(iY[5]),
    .B(iX[23]),
    .Y(_10542_));
 sky130_fd_sc_hd__xnor2_2 _20984_ (.A(_10541_),
    .B(_10542_),
    .Y(_10543_));
 sky130_fd_sc_hd__xnor2_2 _20985_ (.A(_10538_),
    .B(_10543_),
    .Y(_10544_));
 sky130_fd_sc_hd__a21o_2 _20986_ (.A1(_10530_),
    .A2(_10531_),
    .B1(_10544_),
    .X(_10545_));
 sky130_fd_sc_hd__nand3_2 _20987_ (.A(_10530_),
    .B(_10531_),
    .C(_10544_),
    .Y(_10546_));
 sky130_fd_sc_hd__o21ba_2 _20988_ (.A1(_10406_),
    .A2(_10408_),
    .B1_N(_10405_),
    .X(_10547_));
 sky130_fd_sc_hd__o21ba_2 _20989_ (.A1(_10396_),
    .A2(_10398_),
    .B1_N(_10395_),
    .X(_10548_));
 sky130_fd_sc_hd__and4_2 _20990_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[21]),
    .D(iX[22]),
    .X(_10549_));
 sky130_fd_sc_hd__a22oi_2 _20991_ (.A1(iY[7]),
    .A2(iX[21]),
    .B1(iX[22]),
    .B2(iY[6]),
    .Y(_10550_));
 sky130_fd_sc_hd__nor2_2 _20992_ (.A(_10549_),
    .B(_10550_),
    .Y(_10551_));
 sky130_fd_sc_hd__nand2_2 _20993_ (.A(iY[8]),
    .B(iX[20]),
    .Y(_10552_));
 sky130_fd_sc_hd__xnor2_2 _20994_ (.A(_10551_),
    .B(_10552_),
    .Y(_10553_));
 sky130_fd_sc_hd__xnor2_2 _20995_ (.A(_10548_),
    .B(_10553_),
    .Y(_10554_));
 sky130_fd_sc_hd__xnor2_2 _20996_ (.A(_10547_),
    .B(_10554_),
    .Y(_10555_));
 sky130_fd_sc_hd__nand3_2 _20997_ (.A(_10545_),
    .B(_10546_),
    .C(_10555_),
    .Y(_10556_));
 sky130_fd_sc_hd__a21o_2 _20998_ (.A1(_10545_),
    .A2(_10546_),
    .B1(_10555_),
    .X(_10557_));
 sky130_fd_sc_hd__nand2_2 _20999_ (.A(_10556_),
    .B(_10557_),
    .Y(_10558_));
 sky130_fd_sc_hd__nand2_2 _21000_ (.A(_10401_),
    .B(_10412_),
    .Y(_10559_));
 sky130_fd_sc_hd__xnor2_2 _21001_ (.A(_10558_),
    .B(_10559_),
    .Y(_10560_));
 sky130_fd_sc_hd__and2b_2 _21002_ (.A_N(_10430_),
    .B(_10429_),
    .X(_10561_));
 sky130_fd_sc_hd__or2b_2 _21003_ (.A(_10404_),
    .B_N(_10409_),
    .X(_10562_));
 sky130_fd_sc_hd__or2b_2 _21004_ (.A(_10403_),
    .B_N(_10410_),
    .X(_10563_));
 sky130_fd_sc_hd__and4_2 _21005_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[15]),
    .D(iX[16]),
    .X(_10564_));
 sky130_fd_sc_hd__a22oi_2 _21006_ (.A1(iY[13]),
    .A2(iX[15]),
    .B1(iX[16]),
    .B2(iY[12]),
    .Y(_10565_));
 sky130_fd_sc_hd__nor2_2 _21007_ (.A(_10564_),
    .B(_10565_),
    .Y(_10566_));
 sky130_fd_sc_hd__nand2_2 _21008_ (.A(iX[14]),
    .B(iY[14]),
    .Y(_10567_));
 sky130_fd_sc_hd__xnor2_2 _21009_ (.A(_10566_),
    .B(_10567_),
    .Y(_10568_));
 sky130_fd_sc_hd__and4_2 _21010_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[18]),
    .D(iX[19]),
    .X(_10569_));
 sky130_fd_sc_hd__a22oi_2 _21011_ (.A1(iY[10]),
    .A2(iX[18]),
    .B1(iX[19]),
    .B2(iY[9]),
    .Y(_10570_));
 sky130_fd_sc_hd__nor2_2 _21012_ (.A(_10569_),
    .B(_10570_),
    .Y(_10571_));
 sky130_fd_sc_hd__nand2_2 _21013_ (.A(iY[11]),
    .B(iX[17]),
    .Y(_10572_));
 sky130_fd_sc_hd__xnor2_2 _21014_ (.A(_10571_),
    .B(_10572_),
    .Y(_10573_));
 sky130_fd_sc_hd__o21ba_2 _21015_ (.A1(_10426_),
    .A2(_10428_),
    .B1_N(_10425_),
    .X(_10574_));
 sky130_fd_sc_hd__xnor2_2 _21016_ (.A(_10573_),
    .B(_10574_),
    .Y(_10575_));
 sky130_fd_sc_hd__and2_2 _21017_ (.A(_10568_),
    .B(_10575_),
    .X(_10576_));
 sky130_fd_sc_hd__nor2_2 _21018_ (.A(_10568_),
    .B(_10575_),
    .Y(_10577_));
 sky130_fd_sc_hd__or2_2 _21019_ (.A(_10576_),
    .B(_10577_),
    .X(_10578_));
 sky130_fd_sc_hd__a21o_2 _21020_ (.A1(_10562_),
    .A2(_10563_),
    .B1(_10578_),
    .X(_10579_));
 sky130_fd_sc_hd__nand3_2 _21021_ (.A(_10562_),
    .B(_10563_),
    .C(_10578_),
    .Y(_10580_));
 sky130_fd_sc_hd__o211ai_2 _21022_ (.A1(_10561_),
    .A2(_10432_),
    .B1(_10579_),
    .C1(_10580_),
    .Y(_10581_));
 sky130_fd_sc_hd__a211o_2 _21023_ (.A1(_10579_),
    .A2(_10580_),
    .B1(_10561_),
    .C1(_10432_),
    .X(_10582_));
 sky130_fd_sc_hd__and3_2 _21024_ (.A(_10560_),
    .B(_10581_),
    .C(_10582_),
    .X(_10583_));
 sky130_fd_sc_hd__inv_2 _21025_ (.A(_10583_),
    .Y(_10584_));
 sky130_fd_sc_hd__a21o_2 _21026_ (.A1(_10581_),
    .A2(_10582_),
    .B1(_10560_),
    .X(_10585_));
 sky130_fd_sc_hd__o211ai_2 _21027_ (.A1(_10529_),
    .A2(_10441_),
    .B1(_10584_),
    .C1(_10585_),
    .Y(_10586_));
 sky130_fd_sc_hd__a211o_2 _21028_ (.A1(_10584_),
    .A2(_10585_),
    .B1(_10529_),
    .C1(_10441_),
    .X(_10587_));
 sky130_fd_sc_hd__nand2_2 _21029_ (.A(_10586_),
    .B(_10587_),
    .Y(_10588_));
 sky130_fd_sc_hd__a21o_2 _21030_ (.A1(_10461_),
    .A2(_10333_),
    .B1(_10471_),
    .X(_10589_));
 sky130_fd_sc_hd__and4_2 _21031_ (.A(iX[6]),
    .B(iX[7]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_10590_));
 sky130_fd_sc_hd__a22oi_2 _21032_ (.A1(iX[7]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[6]),
    .Y(_10591_));
 sky130_fd_sc_hd__nor2_2 _21033_ (.A(_10590_),
    .B(_10591_),
    .Y(_10592_));
 sky130_fd_sc_hd__nand2_2 _21034_ (.A(iX[5]),
    .B(iY[23]),
    .Y(_10593_));
 sky130_fd_sc_hd__xnor2_2 _21035_ (.A(_10592_),
    .B(_10593_),
    .Y(_10594_));
 sky130_fd_sc_hd__and4_2 _21036_ (.A(iX[9]),
    .B(iX[10]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_10595_));
 sky130_fd_sc_hd__a22oi_2 _21037_ (.A1(iX[10]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[9]),
    .Y(_10596_));
 sky130_fd_sc_hd__nor2_2 _21038_ (.A(_10595_),
    .B(_10596_),
    .Y(_10597_));
 sky130_fd_sc_hd__nand2_2 _21039_ (.A(iX[8]),
    .B(iY[20]),
    .Y(_10598_));
 sky130_fd_sc_hd__xnor2_2 _21040_ (.A(_10597_),
    .B(_10598_),
    .Y(_10599_));
 sky130_fd_sc_hd__o21ba_2 _21041_ (.A1(_10452_),
    .A2(_10454_),
    .B1_N(_10451_),
    .X(_10600_));
 sky130_fd_sc_hd__xnor2_2 _21042_ (.A(_10599_),
    .B(_10600_),
    .Y(_10601_));
 sky130_fd_sc_hd__and2_2 _21043_ (.A(_10594_),
    .B(_10601_),
    .X(_10602_));
 sky130_fd_sc_hd__nor2_2 _21044_ (.A(_10594_),
    .B(_10601_),
    .Y(_10603_));
 sky130_fd_sc_hd__or2_2 _21045_ (.A(_10602_),
    .B(_10603_),
    .X(_10604_));
 sky130_fd_sc_hd__or3_2 _21046_ (.A(_10462_),
    .B(_10465_),
    .C(_10466_),
    .X(_10605_));
 sky130_fd_sc_hd__o21ba_2 _21047_ (.A1(_10421_),
    .A2(_10423_),
    .B1_N(_10420_),
    .X(_10606_));
 sky130_fd_sc_hd__nand4_2 _21048_ (.A(iX[12]),
    .B(iX[13]),
    .C(iY[15]),
    .D(iY[16]),
    .Y(_10607_));
 sky130_fd_sc_hd__a22o_2 _21049_ (.A1(iX[13]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[12]),
    .X(_10608_));
 sky130_fd_sc_hd__and2_2 _21050_ (.A(iX[11]),
    .B(iY[17]),
    .X(_10609_));
 sky130_fd_sc_hd__a21oi_2 _21051_ (.A1(_10607_),
    .A2(_10608_),
    .B1(_10609_),
    .Y(_10610_));
 sky130_fd_sc_hd__and3_2 _21052_ (.A(_10607_),
    .B(_10608_),
    .C(_10609_),
    .X(_10611_));
 sky130_fd_sc_hd__nor2_2 _21053_ (.A(_10610_),
    .B(_10611_),
    .Y(_10612_));
 sky130_fd_sc_hd__xnor2_2 _21054_ (.A(_10606_),
    .B(_10612_),
    .Y(_10613_));
 sky130_fd_sc_hd__o21ai_2 _21055_ (.A1(_10463_),
    .A2(_10465_),
    .B1(_10613_),
    .Y(_10614_));
 sky130_fd_sc_hd__or3_2 _21056_ (.A(_10463_),
    .B(_10465_),
    .C(_10613_),
    .X(_10615_));
 sky130_fd_sc_hd__nand2_2 _21057_ (.A(_10614_),
    .B(_10615_),
    .Y(_10616_));
 sky130_fd_sc_hd__a21oi_2 _21058_ (.A1(_10605_),
    .A2(_10469_),
    .B1(_10616_),
    .Y(_10617_));
 sky130_fd_sc_hd__and3_2 _21059_ (.A(_10605_),
    .B(_10469_),
    .C(_10616_),
    .X(_10618_));
 sky130_fd_sc_hd__or3_2 _21060_ (.A(_10604_),
    .B(_10617_),
    .C(_10618_),
    .X(_10619_));
 sky130_fd_sc_hd__o21ai_2 _21061_ (.A1(_10617_),
    .A2(_10618_),
    .B1(_10604_),
    .Y(_10620_));
 sky130_fd_sc_hd__nand2_2 _21062_ (.A(_10619_),
    .B(_10620_),
    .Y(_10621_));
 sky130_fd_sc_hd__a21oi_2 _21063_ (.A1(_10435_),
    .A2(_10438_),
    .B1(_10621_),
    .Y(_10622_));
 sky130_fd_sc_hd__and3_2 _21064_ (.A(_10435_),
    .B(_10438_),
    .C(_10621_),
    .X(_10623_));
 sky130_fd_sc_hd__a211oi_2 _21065_ (.A1(_10589_),
    .A2(_10474_),
    .B1(_10622_),
    .C1(_10623_),
    .Y(_10624_));
 sky130_fd_sc_hd__o211a_2 _21066_ (.A1(_10622_),
    .A2(_10623_),
    .B1(_10589_),
    .C1(_10474_),
    .X(_10625_));
 sky130_fd_sc_hd__or3_2 _21067_ (.A(_10588_),
    .B(_10624_),
    .C(_10625_),
    .X(_10626_));
 sky130_fd_sc_hd__o21a_2 _21068_ (.A1(_10624_),
    .A2(_10625_),
    .B1(_10588_),
    .X(_10627_));
 sky130_fd_sc_hd__inv_2 _21069_ (.A(_10627_),
    .Y(_10628_));
 sky130_fd_sc_hd__nand2_2 _21070_ (.A(_10626_),
    .B(_10628_),
    .Y(_10629_));
 sky130_fd_sc_hd__a21boi_2 _21071_ (.A1(_10443_),
    .A2(_10444_),
    .B1_N(_10481_),
    .Y(_10630_));
 sky130_fd_sc_hd__xor2_2 _21072_ (.A(_10629_),
    .B(_10630_),
    .X(_10631_));
 sky130_fd_sc_hd__a22o_2 _21073_ (.A1(iX[1]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[0]),
    .X(_10632_));
 sky130_fd_sc_hd__and4_2 _21074_ (.A(iX[0]),
    .B(iX[1]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_10633_));
 sky130_fd_sc_hd__inv_2 _21075_ (.A(_10633_),
    .Y(_10634_));
 sky130_fd_sc_hd__or2b_2 _21076_ (.A(_10488_),
    .B_N(_10493_),
    .X(_10635_));
 sky130_fd_sc_hd__or2b_2 _21077_ (.A(_10487_),
    .B_N(_10494_),
    .X(_10636_));
 sky130_fd_sc_hd__and2b_2 _21078_ (.A_N(_10456_),
    .B(_10455_),
    .X(_10637_));
 sky130_fd_sc_hd__o21ba_2 _21079_ (.A1(_10490_),
    .A2(_10492_),
    .B1_N(_10489_),
    .X(_10638_));
 sky130_fd_sc_hd__o21ba_2 _21080_ (.A1(_10447_),
    .A2(_10449_),
    .B1_N(_10446_),
    .X(_10639_));
 sky130_fd_sc_hd__and4_2 _21081_ (.A(iX[3]),
    .B(iX[4]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_10640_));
 sky130_fd_sc_hd__a22oi_2 _21082_ (.A1(iX[4]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[3]),
    .Y(_10641_));
 sky130_fd_sc_hd__nor2_2 _21083_ (.A(_10640_),
    .B(_10641_),
    .Y(_10642_));
 sky130_fd_sc_hd__nand2_2 _21084_ (.A(iX[2]),
    .B(iY[26]),
    .Y(_10643_));
 sky130_fd_sc_hd__xnor2_2 _21085_ (.A(_10642_),
    .B(_10643_),
    .Y(_10644_));
 sky130_fd_sc_hd__xnor2_2 _21086_ (.A(_10639_),
    .B(_10644_),
    .Y(_10645_));
 sky130_fd_sc_hd__xnor2_2 _21087_ (.A(_10638_),
    .B(_10645_),
    .Y(_10646_));
 sky130_fd_sc_hd__o21a_2 _21088_ (.A1(_10637_),
    .A2(_10458_),
    .B1(_10646_),
    .X(_10647_));
 sky130_fd_sc_hd__nor3_2 _21089_ (.A(_10637_),
    .B(_10458_),
    .C(_10646_),
    .Y(_10648_));
 sky130_fd_sc_hd__a211oi_2 _21090_ (.A1(_10635_),
    .A2(_10636_),
    .B1(_10647_),
    .C1(_10648_),
    .Y(_10649_));
 sky130_fd_sc_hd__o211a_2 _21091_ (.A1(_10647_),
    .A2(_10648_),
    .B1(_10635_),
    .C1(_10636_),
    .X(_10650_));
 sky130_fd_sc_hd__nor2_2 _21092_ (.A(_10496_),
    .B(_10500_),
    .Y(_10651_));
 sky130_fd_sc_hd__or3_2 _21093_ (.A(_10649_),
    .B(_10650_),
    .C(_10651_),
    .X(_10652_));
 sky130_fd_sc_hd__o21ai_2 _21094_ (.A1(_10649_),
    .A2(_10650_),
    .B1(_10651_),
    .Y(_10653_));
 sky130_fd_sc_hd__nand4_2 _21095_ (.A(_10632_),
    .B(_10634_),
    .C(_10652_),
    .D(_10653_),
    .Y(_10654_));
 sky130_fd_sc_hd__a22o_2 _21096_ (.A1(_10632_),
    .A2(_10634_),
    .B1(_10652_),
    .B2(_10653_),
    .X(_10655_));
 sky130_fd_sc_hd__o211a_2 _21097_ (.A1(_10476_),
    .A2(_10479_),
    .B1(_10654_),
    .C1(_10655_),
    .X(_10656_));
 sky130_fd_sc_hd__a211oi_2 _21098_ (.A1(_10654_),
    .A2(_10655_),
    .B1(_10476_),
    .C1(_10479_),
    .Y(_10657_));
 sky130_fd_sc_hd__a211oi_2 _21099_ (.A1(_10504_),
    .A2(_10508_),
    .B1(_10656_),
    .C1(_10657_),
    .Y(_10658_));
 sky130_fd_sc_hd__o211a_2 _21100_ (.A1(_10656_),
    .A2(_10657_),
    .B1(_10504_),
    .C1(_10508_),
    .X(_10659_));
 sky130_fd_sc_hd__nor2_2 _21101_ (.A(_10658_),
    .B(_10659_),
    .Y(_10660_));
 sky130_fd_sc_hd__xnor2_2 _21102_ (.A(_10631_),
    .B(_10660_),
    .Y(_10661_));
 sky130_fd_sc_hd__a21oi_2 _21103_ (.A1(_10484_),
    .A2(_10515_),
    .B1(_10661_),
    .Y(_10662_));
 sky130_fd_sc_hd__and3_2 _21104_ (.A(_10484_),
    .B(_10515_),
    .C(_10661_),
    .X(_10663_));
 sky130_fd_sc_hd__a211oi_2 _21105_ (.A1(_10528_),
    .A2(_10514_),
    .B1(_10662_),
    .C1(_10663_),
    .Y(_10664_));
 sky130_fd_sc_hd__o211a_2 _21106_ (.A1(_10662_),
    .A2(_10663_),
    .B1(_10528_),
    .C1(_10514_),
    .X(_10665_));
 sky130_fd_sc_hd__or2_2 _21107_ (.A(_10664_),
    .B(_10665_),
    .X(_10666_));
 sky130_fd_sc_hd__nand2_2 _21108_ (.A(_10517_),
    .B(_10519_),
    .Y(_10667_));
 sky130_fd_sc_hd__xnor2_2 _21109_ (.A(_10666_),
    .B(_10667_),
    .Y(_10668_));
 sky130_fd_sc_hd__xnor2_2 _21110_ (.A(_10521_),
    .B(_10668_),
    .Y(_10669_));
 sky130_fd_sc_hd__o31a_2 _21111_ (.A1(_10526_),
    .A2(_10380_),
    .A3(_10523_),
    .B1(_10524_),
    .X(_10670_));
 sky130_fd_sc_hd__xnor2_2 _21112_ (.A(_10669_),
    .B(_10670_),
    .Y(_10671_));
 sky130_fd_sc_hd__inv_2 _21113_ (.A(_10671_),
    .Y(oO[28]));
 sky130_fd_sc_hd__and2b_2 _21114_ (.A_N(_10521_),
    .B(_10668_),
    .X(_10672_));
 sky130_fd_sc_hd__o311a_2 _21115_ (.A1(_10526_),
    .A2(_10380_),
    .A3(_10523_),
    .B1(_10524_),
    .C1(_10669_),
    .X(_10673_));
 sky130_fd_sc_hd__and2b_2 _21116_ (.A_N(_10666_),
    .B(_10667_),
    .X(_10674_));
 sky130_fd_sc_hd__and3_2 _21117_ (.A(_10556_),
    .B(_10557_),
    .C(_10559_),
    .X(_10675_));
 sky130_fd_sc_hd__and2b_2 _21118_ (.A_N(_10574_),
    .B(_10573_),
    .X(_10676_));
 sky130_fd_sc_hd__or2b_2 _21119_ (.A(_10548_),
    .B_N(_10553_),
    .X(_10677_));
 sky130_fd_sc_hd__or2b_2 _21120_ (.A(_10547_),
    .B_N(_10554_),
    .X(_10678_));
 sky130_fd_sc_hd__and4_2 _21121_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[16]),
    .D(iX[17]),
    .X(_10679_));
 sky130_fd_sc_hd__a22oi_2 _21122_ (.A1(iY[13]),
    .A2(iX[16]),
    .B1(iX[17]),
    .B2(iY[12]),
    .Y(_10680_));
 sky130_fd_sc_hd__nor2_2 _21123_ (.A(_10679_),
    .B(_10680_),
    .Y(_10681_));
 sky130_fd_sc_hd__nand2_2 _21124_ (.A(iY[14]),
    .B(iX[15]),
    .Y(_10682_));
 sky130_fd_sc_hd__xnor2_2 _21125_ (.A(_10681_),
    .B(_10682_),
    .Y(_10683_));
 sky130_fd_sc_hd__and4_2 _21126_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[19]),
    .D(iX[20]),
    .X(_10684_));
 sky130_fd_sc_hd__a22oi_2 _21127_ (.A1(iY[10]),
    .A2(iX[19]),
    .B1(iX[20]),
    .B2(iY[9]),
    .Y(_10685_));
 sky130_fd_sc_hd__nor2_2 _21128_ (.A(_10684_),
    .B(_10685_),
    .Y(_10686_));
 sky130_fd_sc_hd__nand2_2 _21129_ (.A(iY[11]),
    .B(iX[18]),
    .Y(_10687_));
 sky130_fd_sc_hd__xnor2_2 _21130_ (.A(_10686_),
    .B(_10687_),
    .Y(_10688_));
 sky130_fd_sc_hd__o21ba_2 _21131_ (.A1(_10570_),
    .A2(_10572_),
    .B1_N(_10569_),
    .X(_10689_));
 sky130_fd_sc_hd__xnor2_2 _21132_ (.A(_10688_),
    .B(_10689_),
    .Y(_10690_));
 sky130_fd_sc_hd__and2_2 _21133_ (.A(_10683_),
    .B(_10690_),
    .X(_10691_));
 sky130_fd_sc_hd__nor2_2 _21134_ (.A(_10683_),
    .B(_10690_),
    .Y(_10692_));
 sky130_fd_sc_hd__or2_2 _21135_ (.A(_10691_),
    .B(_10692_),
    .X(_10693_));
 sky130_fd_sc_hd__a21o_2 _21136_ (.A1(_10677_),
    .A2(_10678_),
    .B1(_10693_),
    .X(_10694_));
 sky130_fd_sc_hd__nand3_2 _21137_ (.A(_10677_),
    .B(_10678_),
    .C(_10693_),
    .Y(_10695_));
 sky130_fd_sc_hd__o211ai_2 _21138_ (.A1(_10676_),
    .A2(_10576_),
    .B1(_10694_),
    .C1(_10695_),
    .Y(_10696_));
 sky130_fd_sc_hd__a211o_2 _21139_ (.A1(_10694_),
    .A2(_10695_),
    .B1(_10676_),
    .C1(_10576_),
    .X(_10697_));
 sky130_fd_sc_hd__or2b_2 _21140_ (.A(_10537_),
    .B_N(_10536_),
    .X(_10698_));
 sky130_fd_sc_hd__nand2_2 _21141_ (.A(_10538_),
    .B(_10543_),
    .Y(_10699_));
 sky130_fd_sc_hd__and4_2 _21142_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[28]),
    .D(iX[29]),
    .X(_10700_));
 sky130_fd_sc_hd__a22oi_2 _21143_ (.A1(iY[1]),
    .A2(iX[28]),
    .B1(iX[29]),
    .B2(iY[0]),
    .Y(_10701_));
 sky130_fd_sc_hd__nor2_2 _21144_ (.A(_10700_),
    .B(_10701_),
    .Y(_10702_));
 sky130_fd_sc_hd__nand2_2 _21145_ (.A(iY[2]),
    .B(iX[27]),
    .Y(_10703_));
 sky130_fd_sc_hd__xnor2_2 _21146_ (.A(_10702_),
    .B(_10703_),
    .Y(_10704_));
 sky130_fd_sc_hd__o21ba_2 _21147_ (.A1(_10533_),
    .A2(_10535_),
    .B1_N(_10532_),
    .X(_10705_));
 sky130_fd_sc_hd__xnor2_2 _21148_ (.A(_10704_),
    .B(_10705_),
    .Y(_10706_));
 sky130_fd_sc_hd__and4_2 _21149_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[25]),
    .D(iX[26]),
    .X(_10707_));
 sky130_fd_sc_hd__a22oi_2 _21150_ (.A1(iY[4]),
    .A2(iX[25]),
    .B1(iX[26]),
    .B2(iY[3]),
    .Y(_10708_));
 sky130_fd_sc_hd__nor2_2 _21151_ (.A(_10707_),
    .B(_10708_),
    .Y(_10709_));
 sky130_fd_sc_hd__nand2_2 _21152_ (.A(iY[5]),
    .B(iX[24]),
    .Y(_10710_));
 sky130_fd_sc_hd__xnor2_2 _21153_ (.A(_10709_),
    .B(_10710_),
    .Y(_10711_));
 sky130_fd_sc_hd__xnor2_2 _21154_ (.A(_10706_),
    .B(_10711_),
    .Y(_10712_));
 sky130_fd_sc_hd__a21o_2 _21155_ (.A1(_10698_),
    .A2(_10699_),
    .B1(_10712_),
    .X(_10713_));
 sky130_fd_sc_hd__nand3_2 _21156_ (.A(_10698_),
    .B(_10699_),
    .C(_10712_),
    .Y(_10714_));
 sky130_fd_sc_hd__o21ba_2 _21157_ (.A1(_10550_),
    .A2(_10552_),
    .B1_N(_10549_),
    .X(_10715_));
 sky130_fd_sc_hd__o21ba_2 _21158_ (.A1(_10540_),
    .A2(_10542_),
    .B1_N(_10539_),
    .X(_10716_));
 sky130_fd_sc_hd__and4_2 _21159_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[22]),
    .D(iX[23]),
    .X(_10717_));
 sky130_fd_sc_hd__a22oi_2 _21160_ (.A1(iY[7]),
    .A2(iX[22]),
    .B1(iX[23]),
    .B2(iY[6]),
    .Y(_10718_));
 sky130_fd_sc_hd__nor2_2 _21161_ (.A(_10717_),
    .B(_10718_),
    .Y(_10719_));
 sky130_fd_sc_hd__nand2_2 _21162_ (.A(iY[8]),
    .B(iX[21]),
    .Y(_10720_));
 sky130_fd_sc_hd__xnor2_2 _21163_ (.A(_10719_),
    .B(_10720_),
    .Y(_10721_));
 sky130_fd_sc_hd__xnor2_2 _21164_ (.A(_10716_),
    .B(_10721_),
    .Y(_10722_));
 sky130_fd_sc_hd__xnor2_2 _21165_ (.A(_10715_),
    .B(_10722_),
    .Y(_10723_));
 sky130_fd_sc_hd__nand3_2 _21166_ (.A(_10713_),
    .B(_10714_),
    .C(_10723_),
    .Y(_10724_));
 sky130_fd_sc_hd__a21o_2 _21167_ (.A1(_10713_),
    .A2(_10714_),
    .B1(_10723_),
    .X(_10725_));
 sky130_fd_sc_hd__nand2_2 _21168_ (.A(_10724_),
    .B(_10725_),
    .Y(_10726_));
 sky130_fd_sc_hd__nand2_2 _21169_ (.A(_10545_),
    .B(_10556_),
    .Y(_10727_));
 sky130_fd_sc_hd__xnor2_2 _21170_ (.A(_10726_),
    .B(_10727_),
    .Y(_10728_));
 sky130_fd_sc_hd__a21o_2 _21171_ (.A1(_10696_),
    .A2(_10697_),
    .B1(_10728_),
    .X(_10729_));
 sky130_fd_sc_hd__and3_2 _21172_ (.A(_10728_),
    .B(_10696_),
    .C(_10697_),
    .X(_10730_));
 sky130_fd_sc_hd__inv_2 _21173_ (.A(_10730_),
    .Y(_10731_));
 sky130_fd_sc_hd__o211ai_2 _21174_ (.A1(_10675_),
    .A2(_10583_),
    .B1(_10729_),
    .C1(_10731_),
    .Y(_10732_));
 sky130_fd_sc_hd__a211o_2 _21175_ (.A1(_10729_),
    .A2(_10731_),
    .B1(_10675_),
    .C1(_10583_),
    .X(_10733_));
 sky130_fd_sc_hd__nand2_2 _21176_ (.A(_10732_),
    .B(_10733_),
    .Y(_10734_));
 sky130_fd_sc_hd__inv_2 _21177_ (.A(_10617_),
    .Y(_10735_));
 sky130_fd_sc_hd__and4_2 _21178_ (.A(iX[7]),
    .B(iX[8]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_10736_));
 sky130_fd_sc_hd__a22oi_2 _21179_ (.A1(iX[8]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[7]),
    .Y(_10737_));
 sky130_fd_sc_hd__nor2_2 _21180_ (.A(_10736_),
    .B(_10737_),
    .Y(_10738_));
 sky130_fd_sc_hd__nand2_2 _21181_ (.A(iX[6]),
    .B(iY[23]),
    .Y(_10739_));
 sky130_fd_sc_hd__xnor2_2 _21182_ (.A(_10738_),
    .B(_10739_),
    .Y(_10740_));
 sky130_fd_sc_hd__and4_2 _21183_ (.A(iX[10]),
    .B(iX[11]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_10741_));
 sky130_fd_sc_hd__a22oi_2 _21184_ (.A1(iX[11]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[10]),
    .Y(_10742_));
 sky130_fd_sc_hd__nor2_2 _21185_ (.A(_10741_),
    .B(_10742_),
    .Y(_10743_));
 sky130_fd_sc_hd__nand2_2 _21186_ (.A(iX[9]),
    .B(iY[20]),
    .Y(_10744_));
 sky130_fd_sc_hd__xnor2_2 _21187_ (.A(_10743_),
    .B(_10744_),
    .Y(_10745_));
 sky130_fd_sc_hd__o21ba_2 _21188_ (.A1(_10596_),
    .A2(_10598_),
    .B1_N(_10595_),
    .X(_10746_));
 sky130_fd_sc_hd__xnor2_2 _21189_ (.A(_10745_),
    .B(_10746_),
    .Y(_10747_));
 sky130_fd_sc_hd__and2_2 _21190_ (.A(_10740_),
    .B(_10747_),
    .X(_10748_));
 sky130_fd_sc_hd__nor2_2 _21191_ (.A(_10740_),
    .B(_10747_),
    .Y(_10749_));
 sky130_fd_sc_hd__or2_2 _21192_ (.A(_10748_),
    .B(_10749_),
    .X(_10750_));
 sky130_fd_sc_hd__or3_2 _21193_ (.A(_10606_),
    .B(_10610_),
    .C(_10611_),
    .X(_10751_));
 sky130_fd_sc_hd__and4_2 _21194_ (.A(iX[12]),
    .B(iX[13]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_10752_));
 sky130_fd_sc_hd__o21ba_2 _21195_ (.A1(_10565_),
    .A2(_10567_),
    .B1_N(_10564_),
    .X(_10753_));
 sky130_fd_sc_hd__nand4_2 _21196_ (.A(iX[13]),
    .B(iX[14]),
    .C(iY[15]),
    .D(iY[16]),
    .Y(_10754_));
 sky130_fd_sc_hd__a22o_2 _21197_ (.A1(iX[14]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[13]),
    .X(_10755_));
 sky130_fd_sc_hd__and2_2 _21198_ (.A(iX[12]),
    .B(iY[17]),
    .X(_10756_));
 sky130_fd_sc_hd__a21oi_2 _21199_ (.A1(_10754_),
    .A2(_10755_),
    .B1(_10756_),
    .Y(_10757_));
 sky130_fd_sc_hd__and3_2 _21200_ (.A(_10754_),
    .B(_10755_),
    .C(_10756_),
    .X(_10758_));
 sky130_fd_sc_hd__nor2_2 _21201_ (.A(_10757_),
    .B(_10758_),
    .Y(_10759_));
 sky130_fd_sc_hd__xnor2_2 _21202_ (.A(_10753_),
    .B(_10759_),
    .Y(_10760_));
 sky130_fd_sc_hd__o21ai_2 _21203_ (.A1(_10752_),
    .A2(_10611_),
    .B1(_10760_),
    .Y(_10761_));
 sky130_fd_sc_hd__or3_2 _21204_ (.A(_10752_),
    .B(_10611_),
    .C(_10760_),
    .X(_10762_));
 sky130_fd_sc_hd__nand2_2 _21205_ (.A(_10761_),
    .B(_10762_),
    .Y(_10763_));
 sky130_fd_sc_hd__a21oi_2 _21206_ (.A1(_10751_),
    .A2(_10614_),
    .B1(_10763_),
    .Y(_10764_));
 sky130_fd_sc_hd__and3_2 _21207_ (.A(_10751_),
    .B(_10614_),
    .C(_10763_),
    .X(_10765_));
 sky130_fd_sc_hd__or3_2 _21208_ (.A(_10750_),
    .B(_10764_),
    .C(_10765_),
    .X(_10766_));
 sky130_fd_sc_hd__o21ai_2 _21209_ (.A1(_10764_),
    .A2(_10765_),
    .B1(_10750_),
    .Y(_10767_));
 sky130_fd_sc_hd__nand2_2 _21210_ (.A(_10766_),
    .B(_10767_),
    .Y(_10768_));
 sky130_fd_sc_hd__a21oi_2 _21211_ (.A1(_10579_),
    .A2(_10581_),
    .B1(_10768_),
    .Y(_10769_));
 sky130_fd_sc_hd__and3_2 _21212_ (.A(_10579_),
    .B(_10581_),
    .C(_10768_),
    .X(_10770_));
 sky130_fd_sc_hd__a211oi_2 _21213_ (.A1(_10735_),
    .A2(_10619_),
    .B1(_10769_),
    .C1(_10770_),
    .Y(_10771_));
 sky130_fd_sc_hd__o211a_2 _21214_ (.A1(_10769_),
    .A2(_10770_),
    .B1(_10735_),
    .C1(_10619_),
    .X(_10772_));
 sky130_fd_sc_hd__or3_2 _21215_ (.A(_10734_),
    .B(_10771_),
    .C(_10772_),
    .X(_10773_));
 sky130_fd_sc_hd__inv_2 _21216_ (.A(_10773_),
    .Y(_10774_));
 sky130_fd_sc_hd__o21a_2 _21217_ (.A1(_10771_),
    .A2(_10772_),
    .B1(_10734_),
    .X(_10775_));
 sky130_fd_sc_hd__a211o_2 _21218_ (.A1(_10586_),
    .A2(_10626_),
    .B1(_10774_),
    .C1(_10775_),
    .X(_10776_));
 sky130_fd_sc_hd__inv_2 _21219_ (.A(_10776_),
    .Y(_10777_));
 sky130_fd_sc_hd__o211a_2 _21220_ (.A1(_10774_),
    .A2(_10775_),
    .B1(_10586_),
    .C1(_10626_),
    .X(_10778_));
 sky130_fd_sc_hd__nor2_2 _21221_ (.A(_10777_),
    .B(_10778_),
    .Y(_10779_));
 sky130_fd_sc_hd__and4_2 _21222_ (.A(iX[1]),
    .B(iX[2]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_10780_));
 sky130_fd_sc_hd__a22oi_2 _21223_ (.A1(iX[2]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[1]),
    .Y(_10781_));
 sky130_fd_sc_hd__nor2_2 _21224_ (.A(_10780_),
    .B(_10781_),
    .Y(_10782_));
 sky130_fd_sc_hd__nand2_2 _21225_ (.A(iX[0]),
    .B(iY[29]),
    .Y(_10783_));
 sky130_fd_sc_hd__xnor2_2 _21226_ (.A(_10782_),
    .B(_10783_),
    .Y(_10784_));
 sky130_fd_sc_hd__nand2_2 _21227_ (.A(_10633_),
    .B(_10784_),
    .Y(_10785_));
 sky130_fd_sc_hd__or2_2 _21228_ (.A(_10633_),
    .B(_10784_),
    .X(_10786_));
 sky130_fd_sc_hd__nand2_2 _21229_ (.A(_10785_),
    .B(_10786_),
    .Y(_10787_));
 sky130_fd_sc_hd__or2b_2 _21230_ (.A(_10639_),
    .B_N(_10644_),
    .X(_10788_));
 sky130_fd_sc_hd__or2b_2 _21231_ (.A(_10638_),
    .B_N(_10645_),
    .X(_10789_));
 sky130_fd_sc_hd__and2b_2 _21232_ (.A_N(_10600_),
    .B(_10599_),
    .X(_10790_));
 sky130_fd_sc_hd__o21ba_2 _21233_ (.A1(_10641_),
    .A2(_10643_),
    .B1_N(_10640_),
    .X(_10791_));
 sky130_fd_sc_hd__o21ba_2 _21234_ (.A1(_10591_),
    .A2(_10593_),
    .B1_N(_10590_),
    .X(_10792_));
 sky130_fd_sc_hd__and4_2 _21235_ (.A(iX[4]),
    .B(iX[5]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_10793_));
 sky130_fd_sc_hd__a22oi_2 _21236_ (.A1(iX[5]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[4]),
    .Y(_10794_));
 sky130_fd_sc_hd__nor2_2 _21237_ (.A(_10793_),
    .B(_10794_),
    .Y(_10795_));
 sky130_fd_sc_hd__nand2_2 _21238_ (.A(iX[3]),
    .B(iY[26]),
    .Y(_10796_));
 sky130_fd_sc_hd__xnor2_2 _21239_ (.A(_10795_),
    .B(_10796_),
    .Y(_10797_));
 sky130_fd_sc_hd__xnor2_2 _21240_ (.A(_10792_),
    .B(_10797_),
    .Y(_10798_));
 sky130_fd_sc_hd__xnor2_2 _21241_ (.A(_10791_),
    .B(_10798_),
    .Y(_10799_));
 sky130_fd_sc_hd__o21a_2 _21242_ (.A1(_10790_),
    .A2(_10602_),
    .B1(_10799_),
    .X(_10800_));
 sky130_fd_sc_hd__nor3_2 _21243_ (.A(_10790_),
    .B(_10602_),
    .C(_10799_),
    .Y(_10802_));
 sky130_fd_sc_hd__a211oi_2 _21244_ (.A1(_10788_),
    .A2(_10789_),
    .B1(_10800_),
    .C1(_10802_),
    .Y(_10803_));
 sky130_fd_sc_hd__o211a_2 _21245_ (.A1(_10800_),
    .A2(_10802_),
    .B1(_10788_),
    .C1(_10789_),
    .X(_10804_));
 sky130_fd_sc_hd__nor2_2 _21246_ (.A(_10803_),
    .B(_10804_),
    .Y(_10805_));
 sky130_fd_sc_hd__o21a_2 _21247_ (.A1(_10647_),
    .A2(_10649_),
    .B1(_10805_),
    .X(_10806_));
 sky130_fd_sc_hd__nor3_2 _21248_ (.A(_10647_),
    .B(_10649_),
    .C(_10805_),
    .Y(_10807_));
 sky130_fd_sc_hd__or3_2 _21249_ (.A(_10787_),
    .B(_10806_),
    .C(_10807_),
    .X(_10808_));
 sky130_fd_sc_hd__o21ai_2 _21250_ (.A1(_10806_),
    .A2(_10807_),
    .B1(_10787_),
    .Y(_10809_));
 sky130_fd_sc_hd__o211a_2 _21251_ (.A1(_10622_),
    .A2(_10624_),
    .B1(_10808_),
    .C1(_10809_),
    .X(_10810_));
 sky130_fd_sc_hd__a211oi_2 _21252_ (.A1(_10808_),
    .A2(_10809_),
    .B1(_10622_),
    .C1(_10624_),
    .Y(_10811_));
 sky130_fd_sc_hd__a211oi_2 _21253_ (.A1(_10652_),
    .A2(_10654_),
    .B1(_10810_),
    .C1(_10811_),
    .Y(_10812_));
 sky130_fd_sc_hd__o211a_2 _21254_ (.A1(_10810_),
    .A2(_10811_),
    .B1(_10652_),
    .C1(_10654_),
    .X(_10813_));
 sky130_fd_sc_hd__nor2_2 _21255_ (.A(_10812_),
    .B(_10813_),
    .Y(_10814_));
 sky130_fd_sc_hd__xnor2_2 _21256_ (.A(_10779_),
    .B(_10814_),
    .Y(_10815_));
 sky130_fd_sc_hd__nor2_2 _21257_ (.A(_10629_),
    .B(_10630_),
    .Y(_10816_));
 sky130_fd_sc_hd__a21o_2 _21258_ (.A1(_10631_),
    .A2(_10660_),
    .B1(_10816_),
    .X(_10817_));
 sky130_fd_sc_hd__xnor2_2 _21259_ (.A(_10815_),
    .B(_10817_),
    .Y(_10818_));
 sky130_fd_sc_hd__nor2_2 _21260_ (.A(_10656_),
    .B(_10658_),
    .Y(_10819_));
 sky130_fd_sc_hd__xnor2_2 _21261_ (.A(_10818_),
    .B(_10819_),
    .Y(_10820_));
 sky130_fd_sc_hd__nor2_2 _21262_ (.A(_10662_),
    .B(_10664_),
    .Y(_10821_));
 sky130_fd_sc_hd__xnor2_2 _21263_ (.A(_10820_),
    .B(_10821_),
    .Y(_10823_));
 sky130_fd_sc_hd__nand2_2 _21264_ (.A(_10674_),
    .B(_10823_),
    .Y(_10824_));
 sky130_fd_sc_hd__or2_2 _21265_ (.A(_10674_),
    .B(_10823_),
    .X(_10825_));
 sky130_fd_sc_hd__nand2_2 _21266_ (.A(_10824_),
    .B(_10825_),
    .Y(_10826_));
 sky130_fd_sc_hd__inv_2 _21267_ (.A(_10826_),
    .Y(_10827_));
 sky130_fd_sc_hd__o21a_2 _21268_ (.A1(_10672_),
    .A2(_10673_),
    .B1(_10827_),
    .X(_10828_));
 sky130_fd_sc_hd__nor3_2 _21269_ (.A(_10672_),
    .B(_10673_),
    .C(_10827_),
    .Y(_10829_));
 sky130_fd_sc_hd__or2_2 _21270_ (.A(_10828_),
    .B(_10829_),
    .X(_10830_));
 sky130_fd_sc_hd__inv_2 _21271_ (.A(_10830_),
    .Y(oO[29]));
 sky130_fd_sc_hd__and2b_2 _21272_ (.A_N(_10821_),
    .B(_10820_),
    .X(_10831_));
 sky130_fd_sc_hd__and2b_2 _21273_ (.A_N(_10815_),
    .B(_10817_),
    .X(_10833_));
 sky130_fd_sc_hd__and2b_2 _21274_ (.A_N(_10819_),
    .B(_10818_),
    .X(_10834_));
 sky130_fd_sc_hd__nand2_2 _21275_ (.A(_10779_),
    .B(_10814_),
    .Y(_10835_));
 sky130_fd_sc_hd__and3_2 _21276_ (.A(_10724_),
    .B(_10725_),
    .C(_10727_),
    .X(_10836_));
 sky130_fd_sc_hd__and2b_2 _21277_ (.A_N(_10689_),
    .B(_10688_),
    .X(_10837_));
 sky130_fd_sc_hd__or2b_2 _21278_ (.A(_10716_),
    .B_N(_10721_),
    .X(_10838_));
 sky130_fd_sc_hd__or2b_2 _21279_ (.A(_10715_),
    .B_N(_10722_),
    .X(_10839_));
 sky130_fd_sc_hd__and4_2 _21280_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[17]),
    .D(iX[18]),
    .X(_10840_));
 sky130_fd_sc_hd__a22oi_2 _21281_ (.A1(iY[13]),
    .A2(iX[17]),
    .B1(iX[18]),
    .B2(iY[12]),
    .Y(_10841_));
 sky130_fd_sc_hd__nor2_2 _21282_ (.A(_10840_),
    .B(_10841_),
    .Y(_10842_));
 sky130_fd_sc_hd__nand2_2 _21283_ (.A(iY[14]),
    .B(iX[16]),
    .Y(_10844_));
 sky130_fd_sc_hd__xnor2_2 _21284_ (.A(_10842_),
    .B(_10844_),
    .Y(_10845_));
 sky130_fd_sc_hd__and4_2 _21285_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[20]),
    .D(iX[21]),
    .X(_10846_));
 sky130_fd_sc_hd__a22oi_2 _21286_ (.A1(iY[10]),
    .A2(iX[20]),
    .B1(iX[21]),
    .B2(iY[9]),
    .Y(_10847_));
 sky130_fd_sc_hd__nor2_2 _21287_ (.A(_10846_),
    .B(_10847_),
    .Y(_10848_));
 sky130_fd_sc_hd__nand2_2 _21288_ (.A(iY[11]),
    .B(iX[19]),
    .Y(_10849_));
 sky130_fd_sc_hd__xnor2_2 _21289_ (.A(_10848_),
    .B(_10849_),
    .Y(_10850_));
 sky130_fd_sc_hd__o21ba_2 _21290_ (.A1(_10685_),
    .A2(_10687_),
    .B1_N(_10684_),
    .X(_10851_));
 sky130_fd_sc_hd__xnor2_2 _21291_ (.A(_10850_),
    .B(_10851_),
    .Y(_10852_));
 sky130_fd_sc_hd__and2_2 _21292_ (.A(_10845_),
    .B(_10852_),
    .X(_10853_));
 sky130_fd_sc_hd__nor2_2 _21293_ (.A(_10845_),
    .B(_10852_),
    .Y(_10854_));
 sky130_fd_sc_hd__or2_2 _21294_ (.A(_10853_),
    .B(_10854_),
    .X(_10855_));
 sky130_fd_sc_hd__a21o_2 _21295_ (.A1(_10838_),
    .A2(_10839_),
    .B1(_10855_),
    .X(_10856_));
 sky130_fd_sc_hd__nand3_2 _21296_ (.A(_10838_),
    .B(_10839_),
    .C(_10855_),
    .Y(_10857_));
 sky130_fd_sc_hd__o211ai_2 _21297_ (.A1(_10837_),
    .A2(_10691_),
    .B1(_10856_),
    .C1(_10857_),
    .Y(_10858_));
 sky130_fd_sc_hd__a211o_2 _21298_ (.A1(_10856_),
    .A2(_10857_),
    .B1(_10837_),
    .C1(_10691_),
    .X(_10859_));
 sky130_fd_sc_hd__or2b_2 _21299_ (.A(_10705_),
    .B_N(_10704_),
    .X(_10860_));
 sky130_fd_sc_hd__nand2_2 _21300_ (.A(_10706_),
    .B(_10711_),
    .Y(_10861_));
 sky130_fd_sc_hd__and4_2 _21301_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[29]),
    .D(iX[30]),
    .X(_10862_));
 sky130_fd_sc_hd__a22oi_2 _21302_ (.A1(iY[1]),
    .A2(iX[29]),
    .B1(iX[30]),
    .B2(iY[0]),
    .Y(_10863_));
 sky130_fd_sc_hd__o2bb2a_2 _21303_ (.A1_N(iY[2]),
    .A2_N(iX[28]),
    .B1(_10862_),
    .B2(_10863_),
    .X(_10865_));
 sky130_fd_sc_hd__and4bb_2 _21304_ (.A_N(_10862_),
    .B_N(_10863_),
    .C(iY[2]),
    .D(iX[28]),
    .X(_10866_));
 sky130_fd_sc_hd__nor2_2 _21305_ (.A(_10865_),
    .B(_10866_),
    .Y(_10867_));
 sky130_fd_sc_hd__o21ba_2 _21306_ (.A1(_10701_),
    .A2(_10703_),
    .B1_N(_10700_),
    .X(_10868_));
 sky130_fd_sc_hd__xnor2_2 _21307_ (.A(_10867_),
    .B(_10868_),
    .Y(_10869_));
 sky130_fd_sc_hd__and4_2 _21308_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[26]),
    .D(iX[27]),
    .X(_10870_));
 sky130_fd_sc_hd__a22oi_2 _21309_ (.A1(iY[4]),
    .A2(iX[26]),
    .B1(iX[27]),
    .B2(iY[3]),
    .Y(_10871_));
 sky130_fd_sc_hd__nor2_2 _21310_ (.A(_10870_),
    .B(_10871_),
    .Y(_10872_));
 sky130_fd_sc_hd__nand2_2 _21311_ (.A(iY[5]),
    .B(iX[25]),
    .Y(_10873_));
 sky130_fd_sc_hd__xnor2_2 _21312_ (.A(_10872_),
    .B(_10873_),
    .Y(_10874_));
 sky130_fd_sc_hd__and2_2 _21313_ (.A(_10869_),
    .B(_10874_),
    .X(_10876_));
 sky130_fd_sc_hd__nor2_2 _21314_ (.A(_10869_),
    .B(_10874_),
    .Y(_10877_));
 sky130_fd_sc_hd__or2_2 _21315_ (.A(_10876_),
    .B(_10877_),
    .X(_10878_));
 sky130_fd_sc_hd__a21o_2 _21316_ (.A1(_10860_),
    .A2(_10861_),
    .B1(_10878_),
    .X(_10879_));
 sky130_fd_sc_hd__nand3_2 _21317_ (.A(_10860_),
    .B(_10861_),
    .C(_10878_),
    .Y(_10880_));
 sky130_fd_sc_hd__o21ba_2 _21318_ (.A1(_10718_),
    .A2(_10720_),
    .B1_N(_10717_),
    .X(_10881_));
 sky130_fd_sc_hd__o21ba_2 _21319_ (.A1(_10708_),
    .A2(_10710_),
    .B1_N(_10707_),
    .X(_10882_));
 sky130_fd_sc_hd__and4_2 _21320_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[23]),
    .D(iX[24]),
    .X(_10883_));
 sky130_fd_sc_hd__a22oi_2 _21321_ (.A1(iY[7]),
    .A2(iX[23]),
    .B1(iX[24]),
    .B2(iY[6]),
    .Y(_10884_));
 sky130_fd_sc_hd__nor2_2 _21322_ (.A(_10883_),
    .B(_10884_),
    .Y(_10885_));
 sky130_fd_sc_hd__nand2_2 _21323_ (.A(iY[8]),
    .B(iX[22]),
    .Y(_10887_));
 sky130_fd_sc_hd__xnor2_2 _21324_ (.A(_10885_),
    .B(_10887_),
    .Y(_10888_));
 sky130_fd_sc_hd__xnor2_2 _21325_ (.A(_10882_),
    .B(_10888_),
    .Y(_10889_));
 sky130_fd_sc_hd__xnor2_2 _21326_ (.A(_10881_),
    .B(_10889_),
    .Y(_10890_));
 sky130_fd_sc_hd__nand3_2 _21327_ (.A(_10879_),
    .B(_10880_),
    .C(_10890_),
    .Y(_10891_));
 sky130_fd_sc_hd__a21o_2 _21328_ (.A1(_10879_),
    .A2(_10880_),
    .B1(_10890_),
    .X(_10892_));
 sky130_fd_sc_hd__nand2_2 _21329_ (.A(_10713_),
    .B(_10724_),
    .Y(_10893_));
 sky130_fd_sc_hd__and3_2 _21330_ (.A(_10891_),
    .B(_10892_),
    .C(_10893_),
    .X(_10894_));
 sky130_fd_sc_hd__a21oi_2 _21331_ (.A1(_10891_),
    .A2(_10892_),
    .B1(_10893_),
    .Y(_10895_));
 sky130_fd_sc_hd__nor2_2 _21332_ (.A(_10894_),
    .B(_10895_),
    .Y(_10896_));
 sky130_fd_sc_hd__a21o_2 _21333_ (.A1(_10858_),
    .A2(_10859_),
    .B1(_10896_),
    .X(_10898_));
 sky130_fd_sc_hd__and3_2 _21334_ (.A(_10896_),
    .B(_10858_),
    .C(_10859_),
    .X(_10899_));
 sky130_fd_sc_hd__inv_2 _21335_ (.A(_10899_),
    .Y(_10900_));
 sky130_fd_sc_hd__o211ai_2 _21336_ (.A1(_10836_),
    .A2(_10730_),
    .B1(_10898_),
    .C1(_10900_),
    .Y(_10901_));
 sky130_fd_sc_hd__a211o_2 _21337_ (.A1(_10898_),
    .A2(_10900_),
    .B1(_10836_),
    .C1(_10730_),
    .X(_10902_));
 sky130_fd_sc_hd__nand2_2 _21338_ (.A(_10901_),
    .B(_10902_),
    .Y(_10903_));
 sky130_fd_sc_hd__inv_2 _21339_ (.A(_10764_),
    .Y(_10904_));
 sky130_fd_sc_hd__and4_2 _21340_ (.A(iX[8]),
    .B(iX[9]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_10905_));
 sky130_fd_sc_hd__a22oi_2 _21341_ (.A1(iX[9]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[8]),
    .Y(_10906_));
 sky130_fd_sc_hd__nor2_2 _21342_ (.A(_10905_),
    .B(_10906_),
    .Y(_10907_));
 sky130_fd_sc_hd__nand2_2 _21343_ (.A(iX[7]),
    .B(iY[23]),
    .Y(_10909_));
 sky130_fd_sc_hd__xnor2_2 _21344_ (.A(_10907_),
    .B(_10909_),
    .Y(_10910_));
 sky130_fd_sc_hd__and4_2 _21345_ (.A(iX[11]),
    .B(iX[12]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_10911_));
 sky130_fd_sc_hd__a22oi_2 _21346_ (.A1(iX[12]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[11]),
    .Y(_10912_));
 sky130_fd_sc_hd__nor2_2 _21347_ (.A(_10911_),
    .B(_10912_),
    .Y(_10913_));
 sky130_fd_sc_hd__nand2_2 _21348_ (.A(iX[10]),
    .B(iY[20]),
    .Y(_10914_));
 sky130_fd_sc_hd__xnor2_2 _21349_ (.A(_10913_),
    .B(_10914_),
    .Y(_10915_));
 sky130_fd_sc_hd__o21ba_2 _21350_ (.A1(_10742_),
    .A2(_10744_),
    .B1_N(_10741_),
    .X(_10916_));
 sky130_fd_sc_hd__xnor2_2 _21351_ (.A(_10915_),
    .B(_10916_),
    .Y(_10917_));
 sky130_fd_sc_hd__and2_2 _21352_ (.A(_10910_),
    .B(_10917_),
    .X(_10918_));
 sky130_fd_sc_hd__nor2_2 _21353_ (.A(_10910_),
    .B(_10917_),
    .Y(_10920_));
 sky130_fd_sc_hd__or2_2 _21354_ (.A(_10918_),
    .B(_10920_),
    .X(_10921_));
 sky130_fd_sc_hd__or3_2 _21355_ (.A(_10753_),
    .B(_10757_),
    .C(_10758_),
    .X(_10922_));
 sky130_fd_sc_hd__and4_2 _21356_ (.A(iX[13]),
    .B(iX[14]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_10923_));
 sky130_fd_sc_hd__o21ba_2 _21357_ (.A1(_10680_),
    .A2(_10682_),
    .B1_N(_10679_),
    .X(_10924_));
 sky130_fd_sc_hd__nand4_2 _21358_ (.A(iX[14]),
    .B(iX[15]),
    .C(iY[15]),
    .D(iY[16]),
    .Y(_10925_));
 sky130_fd_sc_hd__a22o_2 _21359_ (.A1(iX[15]),
    .A2(iY[15]),
    .B1(iY[16]),
    .B2(iX[14]),
    .X(_10926_));
 sky130_fd_sc_hd__and2_2 _21360_ (.A(iX[13]),
    .B(iY[17]),
    .X(_10927_));
 sky130_fd_sc_hd__a21oi_2 _21361_ (.A1(_10925_),
    .A2(_10926_),
    .B1(_10927_),
    .Y(_10928_));
 sky130_fd_sc_hd__and3_2 _21362_ (.A(_10925_),
    .B(_10926_),
    .C(_10927_),
    .X(_10929_));
 sky130_fd_sc_hd__nor2_2 _21363_ (.A(_10928_),
    .B(_10929_),
    .Y(_10931_));
 sky130_fd_sc_hd__xnor2_2 _21364_ (.A(_10924_),
    .B(_10931_),
    .Y(_10932_));
 sky130_fd_sc_hd__o21ai_2 _21365_ (.A1(_10923_),
    .A2(_10758_),
    .B1(_10932_),
    .Y(_10933_));
 sky130_fd_sc_hd__or3_2 _21366_ (.A(_10923_),
    .B(_10758_),
    .C(_10932_),
    .X(_10934_));
 sky130_fd_sc_hd__nand2_2 _21367_ (.A(_10933_),
    .B(_10934_),
    .Y(_10935_));
 sky130_fd_sc_hd__a21oi_2 _21368_ (.A1(_10922_),
    .A2(_10761_),
    .B1(_10935_),
    .Y(_10936_));
 sky130_fd_sc_hd__and3_2 _21369_ (.A(_10922_),
    .B(_10761_),
    .C(_10935_),
    .X(_10937_));
 sky130_fd_sc_hd__or3_2 _21370_ (.A(_10921_),
    .B(_10936_),
    .C(_10937_),
    .X(_10938_));
 sky130_fd_sc_hd__o21ai_2 _21371_ (.A1(_10936_),
    .A2(_10937_),
    .B1(_10921_),
    .Y(_10939_));
 sky130_fd_sc_hd__nand2_2 _21372_ (.A(_10938_),
    .B(_10939_),
    .Y(_10940_));
 sky130_fd_sc_hd__a21oi_2 _21373_ (.A1(_10694_),
    .A2(_10696_),
    .B1(_10940_),
    .Y(_10942_));
 sky130_fd_sc_hd__and3_2 _21374_ (.A(_10694_),
    .B(_10696_),
    .C(_10940_),
    .X(_10943_));
 sky130_fd_sc_hd__a211oi_2 _21375_ (.A1(_10904_),
    .A2(_10766_),
    .B1(_10942_),
    .C1(_10943_),
    .Y(_10944_));
 sky130_fd_sc_hd__o211a_2 _21376_ (.A1(_10942_),
    .A2(_10943_),
    .B1(_10904_),
    .C1(_10766_),
    .X(_10945_));
 sky130_fd_sc_hd__or3_2 _21377_ (.A(_10903_),
    .B(_10944_),
    .C(_10945_),
    .X(_10946_));
 sky130_fd_sc_hd__inv_2 _21378_ (.A(_10946_),
    .Y(_10947_));
 sky130_fd_sc_hd__o21a_2 _21379_ (.A1(_10944_),
    .A2(_10945_),
    .B1(_10903_),
    .X(_10948_));
 sky130_fd_sc_hd__a211oi_2 _21380_ (.A1(_10732_),
    .A2(_10773_),
    .B1(_10947_),
    .C1(_10948_),
    .Y(_10949_));
 sky130_fd_sc_hd__o211a_2 _21381_ (.A1(_10947_),
    .A2(_10948_),
    .B1(_10732_),
    .C1(_10773_),
    .X(_10950_));
 sky130_fd_sc_hd__inv_2 _21382_ (.A(_10806_),
    .Y(_10951_));
 sky130_fd_sc_hd__and4_2 _21383_ (.A(iX[2]),
    .B(iX[3]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_10952_));
 sky130_fd_sc_hd__a22o_2 _21384_ (.A1(iX[3]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[2]),
    .X(_10953_));
 sky130_fd_sc_hd__and2b_2 _21385_ (.A_N(_10952_),
    .B(_10953_),
    .X(_10954_));
 sky130_fd_sc_hd__nand2_2 _21386_ (.A(iX[1]),
    .B(iY[29]),
    .Y(_10955_));
 sky130_fd_sc_hd__xnor2_2 _21387_ (.A(_10954_),
    .B(_10955_),
    .Y(_10956_));
 sky130_fd_sc_hd__o21ba_2 _21388_ (.A1(_10781_),
    .A2(_10783_),
    .B1_N(_10780_),
    .X(_10957_));
 sky130_fd_sc_hd__xnor2_2 _21389_ (.A(_10956_),
    .B(_10957_),
    .Y(_10958_));
 sky130_fd_sc_hd__nand3_2 _21390_ (.A(iX[0]),
    .B(iY[30]),
    .C(_10958_),
    .Y(_10959_));
 sky130_fd_sc_hd__a21o_2 _21391_ (.A1(iX[0]),
    .A2(iY[30]),
    .B1(_10958_),
    .X(_10960_));
 sky130_fd_sc_hd__nand2_2 _21392_ (.A(_10959_),
    .B(_10960_),
    .Y(_10961_));
 sky130_fd_sc_hd__or2_2 _21393_ (.A(_10785_),
    .B(_10961_),
    .X(_10963_));
 sky130_fd_sc_hd__nand2_2 _21394_ (.A(_10785_),
    .B(_10961_),
    .Y(_10964_));
 sky130_fd_sc_hd__nand2_2 _21395_ (.A(_10963_),
    .B(_10964_),
    .Y(_10965_));
 sky130_fd_sc_hd__or2b_2 _21396_ (.A(_10792_),
    .B_N(_10797_),
    .X(_10966_));
 sky130_fd_sc_hd__or2b_2 _21397_ (.A(_10791_),
    .B_N(_10798_),
    .X(_10967_));
 sky130_fd_sc_hd__and2b_2 _21398_ (.A_N(_10746_),
    .B(_10745_),
    .X(_10968_));
 sky130_fd_sc_hd__o21ba_2 _21399_ (.A1(_10794_),
    .A2(_10796_),
    .B1_N(_10793_),
    .X(_10969_));
 sky130_fd_sc_hd__o21ba_2 _21400_ (.A1(_10737_),
    .A2(_10739_),
    .B1_N(_10736_),
    .X(_10970_));
 sky130_fd_sc_hd__and4_2 _21401_ (.A(iX[5]),
    .B(iX[6]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_10971_));
 sky130_fd_sc_hd__a22oi_2 _21402_ (.A1(iX[6]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[5]),
    .Y(_10972_));
 sky130_fd_sc_hd__nor2_2 _21403_ (.A(_10971_),
    .B(_10972_),
    .Y(_10974_));
 sky130_fd_sc_hd__nand2_2 _21404_ (.A(iX[4]),
    .B(iY[26]),
    .Y(_10975_));
 sky130_fd_sc_hd__xnor2_2 _21405_ (.A(_10974_),
    .B(_10975_),
    .Y(_10976_));
 sky130_fd_sc_hd__xnor2_2 _21406_ (.A(_10970_),
    .B(_10976_),
    .Y(_10977_));
 sky130_fd_sc_hd__xnor2_2 _21407_ (.A(_10969_),
    .B(_10977_),
    .Y(_10978_));
 sky130_fd_sc_hd__o21a_2 _21408_ (.A1(_10968_),
    .A2(_10748_),
    .B1(_10978_),
    .X(_10979_));
 sky130_fd_sc_hd__nor3_2 _21409_ (.A(_10968_),
    .B(_10748_),
    .C(_10978_),
    .Y(_10980_));
 sky130_fd_sc_hd__a211oi_2 _21410_ (.A1(_10966_),
    .A2(_10967_),
    .B1(_10979_),
    .C1(_10980_),
    .Y(_10981_));
 sky130_fd_sc_hd__o211a_2 _21411_ (.A1(_10979_),
    .A2(_10980_),
    .B1(_10966_),
    .C1(_10967_),
    .X(_10982_));
 sky130_fd_sc_hd__nor2_2 _21412_ (.A(_10981_),
    .B(_10982_),
    .Y(_10983_));
 sky130_fd_sc_hd__o21a_2 _21413_ (.A1(_10800_),
    .A2(_10803_),
    .B1(_10983_),
    .X(_10985_));
 sky130_fd_sc_hd__nor3_2 _21414_ (.A(_10800_),
    .B(_10803_),
    .C(_10983_),
    .Y(_10986_));
 sky130_fd_sc_hd__or3_2 _21415_ (.A(_10965_),
    .B(_10985_),
    .C(_10986_),
    .X(_10987_));
 sky130_fd_sc_hd__o21ai_2 _21416_ (.A1(_10985_),
    .A2(_10986_),
    .B1(_10965_),
    .Y(_10988_));
 sky130_fd_sc_hd__o211a_2 _21417_ (.A1(_10769_),
    .A2(_10771_),
    .B1(_10987_),
    .C1(_10988_),
    .X(_10989_));
 sky130_fd_sc_hd__a211oi_2 _21418_ (.A1(_10987_),
    .A2(_10988_),
    .B1(_10769_),
    .C1(_10771_),
    .Y(_10990_));
 sky130_fd_sc_hd__or2_2 _21419_ (.A(_10989_),
    .B(_10990_),
    .X(_10991_));
 sky130_fd_sc_hd__a21oi_2 _21420_ (.A1(_10951_),
    .A2(_10808_),
    .B1(_10991_),
    .Y(_10992_));
 sky130_fd_sc_hd__and3_2 _21421_ (.A(_10951_),
    .B(_10808_),
    .C(_10991_),
    .X(_10993_));
 sky130_fd_sc_hd__nor4_2 _21422_ (.A(_10949_),
    .B(_10950_),
    .C(_10992_),
    .D(_10993_),
    .Y(_10994_));
 sky130_fd_sc_hd__o22a_2 _21423_ (.A1(_10949_),
    .A2(_10950_),
    .B1(_10992_),
    .B2(_10993_),
    .X(_10996_));
 sky130_fd_sc_hd__a211oi_2 _21424_ (.A1(_10776_),
    .A2(_10835_),
    .B1(_10994_),
    .C1(_10996_),
    .Y(_10997_));
 sky130_fd_sc_hd__o211a_2 _21425_ (.A1(_10994_),
    .A2(_10996_),
    .B1(_10776_),
    .C1(_10835_),
    .X(_10998_));
 sky130_fd_sc_hd__nor2_2 _21426_ (.A(_10997_),
    .B(_10998_),
    .Y(_10999_));
 sky130_fd_sc_hd__nor2_2 _21427_ (.A(_10810_),
    .B(_10812_),
    .Y(_11000_));
 sky130_fd_sc_hd__xnor2_2 _21428_ (.A(_10999_),
    .B(_11000_),
    .Y(_11001_));
 sky130_fd_sc_hd__o21ai_2 _21429_ (.A1(_10833_),
    .A2(_10834_),
    .B1(_11001_),
    .Y(_11002_));
 sky130_fd_sc_hd__or3_2 _21430_ (.A(_10833_),
    .B(_10834_),
    .C(_11001_),
    .X(_11003_));
 sky130_fd_sc_hd__and3_2 _21431_ (.A(_10831_),
    .B(_11002_),
    .C(_11003_),
    .X(_11004_));
 sky130_fd_sc_hd__and2_2 _21432_ (.A(_11002_),
    .B(_11003_),
    .X(_11005_));
 sky130_fd_sc_hd__nor2_2 _21433_ (.A(_10831_),
    .B(_11005_),
    .Y(_11007_));
 sky130_fd_sc_hd__nor2_2 _21434_ (.A(_11004_),
    .B(_11007_),
    .Y(_11008_));
 sky130_fd_sc_hd__inv_2 _21435_ (.A(_10824_),
    .Y(_11009_));
 sky130_fd_sc_hd__nor2_2 _21436_ (.A(_11009_),
    .B(_10828_),
    .Y(_11010_));
 sky130_fd_sc_hd__xnor2_2 _21437_ (.A(_11008_),
    .B(_11010_),
    .Y(oO[30]));
 sky130_fd_sc_hd__o21a_2 _21438_ (.A1(_11009_),
    .A2(_10828_),
    .B1(_11008_),
    .X(_11011_));
 sky130_fd_sc_hd__and2b_2 _21439_ (.A_N(_10851_),
    .B(_10850_),
    .X(_11012_));
 sky130_fd_sc_hd__or2b_2 _21440_ (.A(_10882_),
    .B_N(_10888_),
    .X(_11013_));
 sky130_fd_sc_hd__or2b_2 _21441_ (.A(_10881_),
    .B_N(_10889_),
    .X(_11014_));
 sky130_fd_sc_hd__and4_2 _21442_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[18]),
    .D(iX[19]),
    .X(_11015_));
 sky130_fd_sc_hd__a22oi_2 _21443_ (.A1(iY[13]),
    .A2(iX[18]),
    .B1(iX[19]),
    .B2(iY[12]),
    .Y(_11017_));
 sky130_fd_sc_hd__nor2_2 _21444_ (.A(_11015_),
    .B(_11017_),
    .Y(_11018_));
 sky130_fd_sc_hd__nand2_2 _21445_ (.A(iY[14]),
    .B(iX[17]),
    .Y(_11019_));
 sky130_fd_sc_hd__xnor2_2 _21446_ (.A(_11018_),
    .B(_11019_),
    .Y(_11020_));
 sky130_fd_sc_hd__and4_2 _21447_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[21]),
    .D(iX[22]),
    .X(_11021_));
 sky130_fd_sc_hd__a22oi_2 _21448_ (.A1(iY[10]),
    .A2(iX[21]),
    .B1(iX[22]),
    .B2(iY[9]),
    .Y(_11022_));
 sky130_fd_sc_hd__nor2_2 _21449_ (.A(_11021_),
    .B(_11022_),
    .Y(_11023_));
 sky130_fd_sc_hd__nand2_2 _21450_ (.A(iY[11]),
    .B(iX[20]),
    .Y(_11024_));
 sky130_fd_sc_hd__xnor2_2 _21451_ (.A(_11023_),
    .B(_11024_),
    .Y(_11025_));
 sky130_fd_sc_hd__o21ba_2 _21452_ (.A1(_10847_),
    .A2(_10849_),
    .B1_N(_10846_),
    .X(_11026_));
 sky130_fd_sc_hd__xnor2_2 _21453_ (.A(_11025_),
    .B(_11026_),
    .Y(_11028_));
 sky130_fd_sc_hd__xnor2_2 _21454_ (.A(_11020_),
    .B(_11028_),
    .Y(_11029_));
 sky130_fd_sc_hd__a21o_2 _21455_ (.A1(_11013_),
    .A2(_11014_),
    .B1(_11029_),
    .X(_11030_));
 sky130_fd_sc_hd__nand3_2 _21456_ (.A(_11013_),
    .B(_11014_),
    .C(_11029_),
    .Y(_11031_));
 sky130_fd_sc_hd__o211ai_2 _21457_ (.A1(_11012_),
    .A2(_10853_),
    .B1(_11030_),
    .C1(_11031_),
    .Y(_11032_));
 sky130_fd_sc_hd__a211o_2 _21458_ (.A1(_11030_),
    .A2(_11031_),
    .B1(_11012_),
    .C1(_10853_),
    .X(_11033_));
 sky130_fd_sc_hd__and2b_2 _21459_ (.A_N(_10868_),
    .B(_10867_),
    .X(_11034_));
 sky130_fd_sc_hd__a22oi_2 _21460_ (.A1(iY[1]),
    .A2(iX[30]),
    .B1(iX[31]),
    .B2(iY[0]),
    .Y(_11035_));
 sky130_fd_sc_hd__and4_2 _21461_ (.A(iY[0]),
    .B(iY[1]),
    .C(iX[30]),
    .D(iX[31]),
    .X(_11036_));
 sky130_fd_sc_hd__nor2_2 _21462_ (.A(_11035_),
    .B(_11036_),
    .Y(_11037_));
 sky130_fd_sc_hd__nand2_2 _21463_ (.A(iY[2]),
    .B(iX[29]),
    .Y(_11039_));
 sky130_fd_sc_hd__xnor2_2 _21464_ (.A(_11037_),
    .B(_11039_),
    .Y(_11040_));
 sky130_fd_sc_hd__or2_2 _21465_ (.A(_10862_),
    .B(_10866_),
    .X(_11041_));
 sky130_fd_sc_hd__xnor2_2 _21466_ (.A(_11040_),
    .B(_11041_),
    .Y(_11042_));
 sky130_fd_sc_hd__and4_2 _21467_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[27]),
    .D(iX[28]),
    .X(_11043_));
 sky130_fd_sc_hd__a22oi_2 _21468_ (.A1(iY[4]),
    .A2(iX[27]),
    .B1(iX[28]),
    .B2(iY[3]),
    .Y(_11044_));
 sky130_fd_sc_hd__nand2_2 _21469_ (.A(iY[5]),
    .B(iX[26]),
    .Y(_11045_));
 sky130_fd_sc_hd__o21a_2 _21470_ (.A1(_11043_),
    .A2(_11044_),
    .B1(_11045_),
    .X(_11046_));
 sky130_fd_sc_hd__nor3_2 _21471_ (.A(_11043_),
    .B(_11044_),
    .C(_11045_),
    .Y(_11047_));
 sky130_fd_sc_hd__nor2_2 _21472_ (.A(_11046_),
    .B(_11047_),
    .Y(_11048_));
 sky130_fd_sc_hd__xnor2_2 _21473_ (.A(_11042_),
    .B(_11048_),
    .Y(_11050_));
 sky130_fd_sc_hd__o21ai_2 _21474_ (.A1(_11034_),
    .A2(_10876_),
    .B1(_11050_),
    .Y(_11051_));
 sky130_fd_sc_hd__or3_2 _21475_ (.A(_11034_),
    .B(_10876_),
    .C(_11050_),
    .X(_11052_));
 sky130_fd_sc_hd__o21ba_2 _21476_ (.A1(_10884_),
    .A2(_10887_),
    .B1_N(_10883_),
    .X(_11053_));
 sky130_fd_sc_hd__o21ba_2 _21477_ (.A1(_10871_),
    .A2(_10873_),
    .B1_N(_10870_),
    .X(_11054_));
 sky130_fd_sc_hd__and4_2 _21478_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[24]),
    .D(iX[25]),
    .X(_11055_));
 sky130_fd_sc_hd__a22oi_2 _21479_ (.A1(iY[7]),
    .A2(iX[24]),
    .B1(iX[25]),
    .B2(iY[6]),
    .Y(_11056_));
 sky130_fd_sc_hd__nor2_2 _21480_ (.A(_11055_),
    .B(_11056_),
    .Y(_11057_));
 sky130_fd_sc_hd__a21oi_2 _21481_ (.A1(iY[8]),
    .A2(iX[23]),
    .B1(_11057_),
    .Y(_11058_));
 sky130_fd_sc_hd__and3_2 _21482_ (.A(iY[8]),
    .B(iX[23]),
    .C(_11057_),
    .X(_11059_));
 sky130_fd_sc_hd__nor2_2 _21483_ (.A(_11058_),
    .B(_11059_),
    .Y(_11061_));
 sky130_fd_sc_hd__xnor2_2 _21484_ (.A(_11054_),
    .B(_11061_),
    .Y(_11062_));
 sky130_fd_sc_hd__xnor2_2 _21485_ (.A(_11053_),
    .B(_11062_),
    .Y(_11063_));
 sky130_fd_sc_hd__nand3_2 _21486_ (.A(_11051_),
    .B(_11052_),
    .C(_11063_),
    .Y(_11064_));
 sky130_fd_sc_hd__a21o_2 _21487_ (.A1(_11051_),
    .A2(_11052_),
    .B1(_11063_),
    .X(_11065_));
 sky130_fd_sc_hd__nand2_2 _21488_ (.A(_10879_),
    .B(_10891_),
    .Y(_11066_));
 sky130_fd_sc_hd__and3_2 _21489_ (.A(_11064_),
    .B(_11065_),
    .C(_11066_),
    .X(_11067_));
 sky130_fd_sc_hd__a21oi_2 _21490_ (.A1(_11064_),
    .A2(_11065_),
    .B1(_11066_),
    .Y(_11068_));
 sky130_fd_sc_hd__nor2_2 _21491_ (.A(_11067_),
    .B(_11068_),
    .Y(_11069_));
 sky130_fd_sc_hd__a21o_2 _21492_ (.A1(_11032_),
    .A2(_11033_),
    .B1(_11069_),
    .X(_11070_));
 sky130_fd_sc_hd__and3_2 _21493_ (.A(_11069_),
    .B(_11032_),
    .C(_11033_),
    .X(_11072_));
 sky130_fd_sc_hd__inv_2 _21494_ (.A(_11072_),
    .Y(_11073_));
 sky130_fd_sc_hd__o211a_2 _21495_ (.A1(_10894_),
    .A2(_10899_),
    .B1(_11070_),
    .C1(_11073_),
    .X(_11074_));
 sky130_fd_sc_hd__a211oi_2 _21496_ (.A1(_11070_),
    .A2(_11073_),
    .B1(_10894_),
    .C1(_10899_),
    .Y(_11075_));
 sky130_fd_sc_hd__inv_2 _21497_ (.A(_10936_),
    .Y(_11076_));
 sky130_fd_sc_hd__and4_2 _21498_ (.A(iX[9]),
    .B(iX[10]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_11077_));
 sky130_fd_sc_hd__a22oi_2 _21499_ (.A1(iX[10]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[9]),
    .Y(_11078_));
 sky130_fd_sc_hd__nor2_2 _21500_ (.A(_11077_),
    .B(_11078_),
    .Y(_11079_));
 sky130_fd_sc_hd__nand2_2 _21501_ (.A(iX[8]),
    .B(iY[23]),
    .Y(_11080_));
 sky130_fd_sc_hd__xnor2_2 _21502_ (.A(_11079_),
    .B(_11080_),
    .Y(_11081_));
 sky130_fd_sc_hd__and4_2 _21503_ (.A(iX[12]),
    .B(iX[13]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_11083_));
 sky130_fd_sc_hd__a22oi_2 _21504_ (.A1(iX[13]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[12]),
    .Y(_11084_));
 sky130_fd_sc_hd__nor2_2 _21505_ (.A(_11083_),
    .B(_11084_),
    .Y(_11085_));
 sky130_fd_sc_hd__nand2_2 _21506_ (.A(iX[11]),
    .B(iY[20]),
    .Y(_11086_));
 sky130_fd_sc_hd__xnor2_2 _21507_ (.A(_11085_),
    .B(_11086_),
    .Y(_11087_));
 sky130_fd_sc_hd__o21ba_2 _21508_ (.A1(_10912_),
    .A2(_10914_),
    .B1_N(_10911_),
    .X(_11088_));
 sky130_fd_sc_hd__xnor2_2 _21509_ (.A(_11087_),
    .B(_11088_),
    .Y(_11089_));
 sky130_fd_sc_hd__and2_2 _21510_ (.A(_11081_),
    .B(_11089_),
    .X(_11090_));
 sky130_fd_sc_hd__nor2_2 _21511_ (.A(_11081_),
    .B(_11089_),
    .Y(_11091_));
 sky130_fd_sc_hd__or2_2 _21512_ (.A(_11090_),
    .B(_11091_),
    .X(_11092_));
 sky130_fd_sc_hd__or3_2 _21513_ (.A(_10924_),
    .B(_10928_),
    .C(_10929_),
    .X(_11094_));
 sky130_fd_sc_hd__and4_2 _21514_ (.A(iX[14]),
    .B(iX[15]),
    .C(iY[15]),
    .D(iY[16]),
    .X(_11095_));
 sky130_fd_sc_hd__o21ba_2 _21515_ (.A1(_10841_),
    .A2(_10844_),
    .B1_N(_10840_),
    .X(_11096_));
 sky130_fd_sc_hd__nand4_2 _21516_ (.A(iX[15]),
    .B(iY[15]),
    .C(iX[16]),
    .D(iY[16]),
    .Y(_11097_));
 sky130_fd_sc_hd__a22o_2 _21517_ (.A1(iY[15]),
    .A2(iX[16]),
    .B1(iY[16]),
    .B2(iX[15]),
    .X(_11098_));
 sky130_fd_sc_hd__and2_2 _21518_ (.A(iX[14]),
    .B(iY[17]),
    .X(_11099_));
 sky130_fd_sc_hd__a21oi_2 _21519_ (.A1(_11097_),
    .A2(_11098_),
    .B1(_11099_),
    .Y(_11100_));
 sky130_fd_sc_hd__and3_2 _21520_ (.A(_11097_),
    .B(_11098_),
    .C(_11099_),
    .X(_11101_));
 sky130_fd_sc_hd__nor2_2 _21521_ (.A(_11100_),
    .B(_11101_),
    .Y(_11102_));
 sky130_fd_sc_hd__xnor2_2 _21522_ (.A(_11096_),
    .B(_11102_),
    .Y(_11103_));
 sky130_fd_sc_hd__o21ai_2 _21523_ (.A1(_11095_),
    .A2(_10929_),
    .B1(_11103_),
    .Y(_11104_));
 sky130_fd_sc_hd__or3_2 _21524_ (.A(_11095_),
    .B(_10929_),
    .C(_11103_),
    .X(_11105_));
 sky130_fd_sc_hd__nand2_2 _21525_ (.A(_11104_),
    .B(_11105_),
    .Y(_11106_));
 sky130_fd_sc_hd__a21oi_2 _21526_ (.A1(_11094_),
    .A2(_10933_),
    .B1(_11106_),
    .Y(_11107_));
 sky130_fd_sc_hd__and3_2 _21527_ (.A(_11094_),
    .B(_10933_),
    .C(_11106_),
    .X(_11108_));
 sky130_fd_sc_hd__nor3_2 _21528_ (.A(_11092_),
    .B(_11107_),
    .C(_11108_),
    .Y(_11109_));
 sky130_fd_sc_hd__o21a_2 _21529_ (.A1(_11107_),
    .A2(_11108_),
    .B1(_11092_),
    .X(_11110_));
 sky130_fd_sc_hd__a211oi_2 _21530_ (.A1(_10856_),
    .A2(_10858_),
    .B1(_11109_),
    .C1(_11110_),
    .Y(_11111_));
 sky130_fd_sc_hd__o211a_2 _21531_ (.A1(_11109_),
    .A2(_11110_),
    .B1(_10856_),
    .C1(_10858_),
    .X(_11112_));
 sky130_fd_sc_hd__a211oi_2 _21532_ (.A1(_11076_),
    .A2(_10938_),
    .B1(_11111_),
    .C1(_11112_),
    .Y(_11113_));
 sky130_fd_sc_hd__o211a_2 _21533_ (.A1(_11111_),
    .A2(_11112_),
    .B1(_11076_),
    .C1(_10938_),
    .X(_11115_));
 sky130_fd_sc_hd__nor4_2 _21534_ (.A(_11074_),
    .B(_11075_),
    .C(_11113_),
    .D(_11115_),
    .Y(_11116_));
 sky130_fd_sc_hd__o22a_2 _21535_ (.A1(_11074_),
    .A2(_11075_),
    .B1(_11113_),
    .B2(_11115_),
    .X(_11117_));
 sky130_fd_sc_hd__a211o_2 _21536_ (.A1(_10901_),
    .A2(_10946_),
    .B1(_11116_),
    .C1(_11117_),
    .X(_11118_));
 sky130_fd_sc_hd__o211ai_2 _21537_ (.A1(_11116_),
    .A2(_11117_),
    .B1(_10901_),
    .C1(_10946_),
    .Y(_11119_));
 sky130_fd_sc_hd__inv_2 _21538_ (.A(_10987_),
    .Y(_11120_));
 sky130_fd_sc_hd__or2b_2 _21539_ (.A(_10957_),
    .B_N(_10956_),
    .X(_11121_));
 sky130_fd_sc_hd__and4_2 _21540_ (.A(iX[3]),
    .B(iX[4]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_11122_));
 sky130_fd_sc_hd__a22oi_2 _21541_ (.A1(iX[4]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[3]),
    .Y(_11123_));
 sky130_fd_sc_hd__nor2_2 _21542_ (.A(_11122_),
    .B(_11123_),
    .Y(_11124_));
 sky130_fd_sc_hd__nand2_2 _21543_ (.A(iX[2]),
    .B(iY[29]),
    .Y(_11126_));
 sky130_fd_sc_hd__xnor2_2 _21544_ (.A(_11124_),
    .B(_11126_),
    .Y(_11127_));
 sky130_fd_sc_hd__a31o_2 _21545_ (.A1(iX[1]),
    .A2(iY[29]),
    .A3(_10953_),
    .B1(_10952_),
    .X(_11128_));
 sky130_fd_sc_hd__and2_2 _21546_ (.A(_11127_),
    .B(_11128_),
    .X(_11129_));
 sky130_fd_sc_hd__nor2_2 _21547_ (.A(_11127_),
    .B(_11128_),
    .Y(_11130_));
 sky130_fd_sc_hd__nor2_2 _21548_ (.A(_11129_),
    .B(_11130_),
    .Y(_11131_));
 sky130_fd_sc_hd__and2_2 _21549_ (.A(iX[1]),
    .B(iY[30]),
    .X(_11132_));
 sky130_fd_sc_hd__nor2_2 _21550_ (.A(_11131_),
    .B(_11132_),
    .Y(_11133_));
 sky130_fd_sc_hd__and2_2 _21551_ (.A(_11131_),
    .B(_11132_),
    .X(_11134_));
 sky130_fd_sc_hd__or2_2 _21552_ (.A(_11133_),
    .B(_11134_),
    .X(_11135_));
 sky130_fd_sc_hd__a21oi_2 _21553_ (.A1(_11121_),
    .A2(_10959_),
    .B1(_11135_),
    .Y(_11137_));
 sky130_fd_sc_hd__and3_2 _21554_ (.A(_11121_),
    .B(_10959_),
    .C(_11135_),
    .X(_11138_));
 sky130_fd_sc_hd__nor2_2 _21555_ (.A(_11137_),
    .B(_11138_),
    .Y(_11139_));
 sky130_fd_sc_hd__nand2_2 _21556_ (.A(iX[0]),
    .B(iY[31]),
    .Y(_11140_));
 sky130_fd_sc_hd__xnor2_2 _21557_ (.A(_11139_),
    .B(_11140_),
    .Y(_11141_));
 sky130_fd_sc_hd__or2b_2 _21558_ (.A(_10970_),
    .B_N(_10976_),
    .X(_11142_));
 sky130_fd_sc_hd__or2b_2 _21559_ (.A(_10969_),
    .B_N(_10977_),
    .X(_11143_));
 sky130_fd_sc_hd__and2b_2 _21560_ (.A_N(_10916_),
    .B(_10915_),
    .X(_11144_));
 sky130_fd_sc_hd__o21ba_2 _21561_ (.A1(_10972_),
    .A2(_10975_),
    .B1_N(_10971_),
    .X(_11145_));
 sky130_fd_sc_hd__o21ba_2 _21562_ (.A1(_10906_),
    .A2(_10909_),
    .B1_N(_10905_),
    .X(_11146_));
 sky130_fd_sc_hd__and4_2 _21563_ (.A(iX[6]),
    .B(iX[7]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_11148_));
 sky130_fd_sc_hd__a22oi_2 _21564_ (.A1(iX[7]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[6]),
    .Y(_11149_));
 sky130_fd_sc_hd__nor2_2 _21565_ (.A(_11148_),
    .B(_11149_),
    .Y(_11150_));
 sky130_fd_sc_hd__nand2_2 _21566_ (.A(iX[5]),
    .B(iY[26]),
    .Y(_11151_));
 sky130_fd_sc_hd__xnor2_2 _21567_ (.A(_11150_),
    .B(_11151_),
    .Y(_11152_));
 sky130_fd_sc_hd__xnor2_2 _21568_ (.A(_11146_),
    .B(_11152_),
    .Y(_11153_));
 sky130_fd_sc_hd__xnor2_2 _21569_ (.A(_11145_),
    .B(_11153_),
    .Y(_11154_));
 sky130_fd_sc_hd__o21a_2 _21570_ (.A1(_11144_),
    .A2(_10918_),
    .B1(_11154_),
    .X(_11155_));
 sky130_fd_sc_hd__nor3_2 _21571_ (.A(_11144_),
    .B(_10918_),
    .C(_11154_),
    .Y(_11156_));
 sky130_fd_sc_hd__a211oi_2 _21572_ (.A1(_11142_),
    .A2(_11143_),
    .B1(_11155_),
    .C1(_11156_),
    .Y(_11157_));
 sky130_fd_sc_hd__o211a_2 _21573_ (.A1(_11155_),
    .A2(_11156_),
    .B1(_11142_),
    .C1(_11143_),
    .X(_11159_));
 sky130_fd_sc_hd__nor2_2 _21574_ (.A(_10979_),
    .B(_10981_),
    .Y(_11160_));
 sky130_fd_sc_hd__or3_2 _21575_ (.A(_11157_),
    .B(_11159_),
    .C(_11160_),
    .X(_11161_));
 sky130_fd_sc_hd__o21ai_2 _21576_ (.A1(_11157_),
    .A2(_11159_),
    .B1(_11160_),
    .Y(_11162_));
 sky130_fd_sc_hd__and3_2 _21577_ (.A(_11141_),
    .B(_11161_),
    .C(_11162_),
    .X(_11163_));
 sky130_fd_sc_hd__a21oi_2 _21578_ (.A1(_11161_),
    .A2(_11162_),
    .B1(_11141_),
    .Y(_11164_));
 sky130_fd_sc_hd__nor2_2 _21579_ (.A(_11163_),
    .B(_11164_),
    .Y(_11165_));
 sky130_fd_sc_hd__o21ai_2 _21580_ (.A1(_10942_),
    .A2(_10944_),
    .B1(_11165_),
    .Y(_11166_));
 sky130_fd_sc_hd__or3_2 _21581_ (.A(_10942_),
    .B(_10944_),
    .C(_11165_),
    .X(_11167_));
 sky130_fd_sc_hd__o211ai_2 _21582_ (.A1(_10985_),
    .A2(_11120_),
    .B1(_11166_),
    .C1(_11167_),
    .Y(_11168_));
 sky130_fd_sc_hd__a211o_2 _21583_ (.A1(_11166_),
    .A2(_11167_),
    .B1(_10985_),
    .C1(_11120_),
    .X(_11170_));
 sky130_fd_sc_hd__nand4_2 _21584_ (.A(_11118_),
    .B(_11119_),
    .C(_11168_),
    .D(_11170_),
    .Y(_11171_));
 sky130_fd_sc_hd__a22o_2 _21585_ (.A1(_11118_),
    .A2(_11119_),
    .B1(_11168_),
    .B2(_11170_),
    .X(_11172_));
 sky130_fd_sc_hd__o211ai_2 _21586_ (.A1(_10949_),
    .A2(_10994_),
    .B1(_11171_),
    .C1(_11172_),
    .Y(_11173_));
 sky130_fd_sc_hd__a211o_2 _21587_ (.A1(_11171_),
    .A2(_11172_),
    .B1(_10949_),
    .C1(_10994_),
    .X(_11174_));
 sky130_fd_sc_hd__o211ai_2 _21588_ (.A1(_10989_),
    .A2(_10992_),
    .B1(_11173_),
    .C1(_11174_),
    .Y(_11175_));
 sky130_fd_sc_hd__a211o_2 _21589_ (.A1(_11173_),
    .A2(_11174_),
    .B1(_10989_),
    .C1(_10992_),
    .X(_11176_));
 sky130_fd_sc_hd__nand2_2 _21590_ (.A(_11175_),
    .B(_11176_),
    .Y(_11177_));
 sky130_fd_sc_hd__o21ba_2 _21591_ (.A1(_10998_),
    .A2(_11000_),
    .B1_N(_10997_),
    .X(_11178_));
 sky130_fd_sc_hd__xnor2_2 _21592_ (.A(_11177_),
    .B(_11178_),
    .Y(_11179_));
 sky130_fd_sc_hd__nor2_2 _21593_ (.A(_10963_),
    .B(_11179_),
    .Y(_11181_));
 sky130_fd_sc_hd__and2_2 _21594_ (.A(_10963_),
    .B(_11179_),
    .X(_11182_));
 sky130_fd_sc_hd__nor2_2 _21595_ (.A(_11181_),
    .B(_11182_),
    .Y(_11183_));
 sky130_fd_sc_hd__xnor2_2 _21596_ (.A(_11002_),
    .B(_11183_),
    .Y(_11184_));
 sky130_fd_sc_hd__o21ai_2 _21597_ (.A1(_11004_),
    .A2(_11011_),
    .B1(_11184_),
    .Y(_11185_));
 sky130_fd_sc_hd__or3_2 _21598_ (.A(_11004_),
    .B(_11011_),
    .C(_11184_),
    .X(_11186_));
 sky130_fd_sc_hd__and2_2 _21599_ (.A(_11185_),
    .B(_11186_),
    .X(_11187_));
 sky130_fd_sc_hd__buf_1 _21600_ (.A(_11187_),
    .X(oO[31]));
 sky130_fd_sc_hd__or2b_2 _21601_ (.A(_11002_),
    .B_N(_11183_),
    .X(_11188_));
 sky130_fd_sc_hd__nor2_2 _21602_ (.A(_11177_),
    .B(_11178_),
    .Y(_11189_));
 sky130_fd_sc_hd__a31o_2 _21603_ (.A1(iX[0]),
    .A2(iY[31]),
    .A3(_11139_),
    .B1(_11137_),
    .X(_11191_));
 sky130_fd_sc_hd__nand2_2 _21604_ (.A(_11166_),
    .B(_11168_),
    .Y(_11192_));
 sky130_fd_sc_hd__or2b_2 _21605_ (.A(_11146_),
    .B_N(_11152_),
    .X(_11193_));
 sky130_fd_sc_hd__or2b_2 _21606_ (.A(_11145_),
    .B_N(_11153_),
    .X(_11194_));
 sky130_fd_sc_hd__nand2_2 _21607_ (.A(_11193_),
    .B(_11194_),
    .Y(_11195_));
 sky130_fd_sc_hd__and2b_2 _21608_ (.A_N(_11088_),
    .B(_11087_),
    .X(_11196_));
 sky130_fd_sc_hd__o21ba_2 _21609_ (.A1(_11149_),
    .A2(_11151_),
    .B1_N(_11148_),
    .X(_11197_));
 sky130_fd_sc_hd__o21ba_2 _21610_ (.A1(_11078_),
    .A2(_11080_),
    .B1_N(_11077_),
    .X(_11198_));
 sky130_fd_sc_hd__nand2_2 _21611_ (.A(iX[6]),
    .B(iY[26]),
    .Y(_11199_));
 sky130_fd_sc_hd__and4_2 _21612_ (.A(iX[7]),
    .B(iX[8]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_11200_));
 sky130_fd_sc_hd__a22oi_2 _21613_ (.A1(iX[8]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[7]),
    .Y(_11202_));
 sky130_fd_sc_hd__nor2_2 _21614_ (.A(_11200_),
    .B(_11202_),
    .Y(_11203_));
 sky130_fd_sc_hd__xnor2_2 _21615_ (.A(_11199_),
    .B(_11203_),
    .Y(_11204_));
 sky130_fd_sc_hd__xnor2_2 _21616_ (.A(_11198_),
    .B(_11204_),
    .Y(_11205_));
 sky130_fd_sc_hd__xnor2_2 _21617_ (.A(_11197_),
    .B(_11205_),
    .Y(_11206_));
 sky130_fd_sc_hd__o21a_2 _21618_ (.A1(_11196_),
    .A2(_11090_),
    .B1(_11206_),
    .X(_11207_));
 sky130_fd_sc_hd__nor3_2 _21619_ (.A(_11196_),
    .B(_11090_),
    .C(_11206_),
    .Y(_11208_));
 sky130_fd_sc_hd__or2_2 _21620_ (.A(_11207_),
    .B(_11208_),
    .X(_11209_));
 sky130_fd_sc_hd__xnor2_2 _21621_ (.A(_11195_),
    .B(_11209_),
    .Y(_11210_));
 sky130_fd_sc_hd__o21ai_2 _21622_ (.A1(_11155_),
    .A2(_11157_),
    .B1(_11210_),
    .Y(_11211_));
 sky130_fd_sc_hd__or3_2 _21623_ (.A(_11155_),
    .B(_11157_),
    .C(_11210_),
    .X(_11213_));
 sky130_fd_sc_hd__nand2_2 _21624_ (.A(iX[1]),
    .B(iY[31]),
    .Y(_11214_));
 sky130_fd_sc_hd__nand2_2 _21625_ (.A(iX[3]),
    .B(iY[29]),
    .Y(_11215_));
 sky130_fd_sc_hd__and4_2 _21626_ (.A(iX[4]),
    .B(iX[5]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_11216_));
 sky130_fd_sc_hd__a22oi_2 _21627_ (.A1(iX[5]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[4]),
    .Y(_11217_));
 sky130_fd_sc_hd__nor2_2 _21628_ (.A(_11216_),
    .B(_11217_),
    .Y(_11218_));
 sky130_fd_sc_hd__xnor2_2 _21629_ (.A(_11215_),
    .B(_11218_),
    .Y(_11219_));
 sky130_fd_sc_hd__o21ba_2 _21630_ (.A1(_11123_),
    .A2(_11126_),
    .B1_N(_11122_),
    .X(_11220_));
 sky130_fd_sc_hd__xnor2_2 _21631_ (.A(_11219_),
    .B(_11220_),
    .Y(_11221_));
 sky130_fd_sc_hd__nand3_2 _21632_ (.A(iX[2]),
    .B(iY[30]),
    .C(_11221_),
    .Y(_11222_));
 sky130_fd_sc_hd__a21o_2 _21633_ (.A1(iX[2]),
    .A2(iY[30]),
    .B1(_11221_),
    .X(_11224_));
 sky130_fd_sc_hd__and2_2 _21634_ (.A(_11222_),
    .B(_11224_),
    .X(_11225_));
 sky130_fd_sc_hd__o21a_2 _21635_ (.A1(_11129_),
    .A2(_11134_),
    .B1(_11225_),
    .X(_11226_));
 sky130_fd_sc_hd__nor3_2 _21636_ (.A(_11129_),
    .B(_11134_),
    .C(_11225_),
    .Y(_11227_));
 sky130_fd_sc_hd__nor2_2 _21637_ (.A(_11226_),
    .B(_11227_),
    .Y(_11228_));
 sky130_fd_sc_hd__xnor2_2 _21638_ (.A(_11214_),
    .B(_11228_),
    .Y(_11229_));
 sky130_fd_sc_hd__and3_2 _21639_ (.A(_11211_),
    .B(_11213_),
    .C(_11229_),
    .X(_11230_));
 sky130_fd_sc_hd__a21oi_2 _21640_ (.A1(_11211_),
    .A2(_11213_),
    .B1(_11229_),
    .Y(_11231_));
 sky130_fd_sc_hd__nor2_2 _21641_ (.A(_11230_),
    .B(_11231_),
    .Y(_11232_));
 sky130_fd_sc_hd__o21ai_2 _21642_ (.A1(_11111_),
    .A2(_11113_),
    .B1(_11232_),
    .Y(_11233_));
 sky130_fd_sc_hd__or3_2 _21643_ (.A(_11111_),
    .B(_11113_),
    .C(_11232_),
    .X(_11235_));
 sky130_fd_sc_hd__nand2_2 _21644_ (.A(_11233_),
    .B(_11235_),
    .Y(_11236_));
 sky130_fd_sc_hd__a21bo_2 _21645_ (.A1(_11141_),
    .A2(_11162_),
    .B1_N(_11161_),
    .X(_11237_));
 sky130_fd_sc_hd__xnor2_2 _21646_ (.A(_11236_),
    .B(_11237_),
    .Y(_11238_));
 sky130_fd_sc_hd__nand2_2 _21647_ (.A(_11030_),
    .B(_11032_),
    .Y(_11239_));
 sky130_fd_sc_hd__or3_2 _21648_ (.A(_11096_),
    .B(_11100_),
    .C(_11101_),
    .X(_11240_));
 sky130_fd_sc_hd__and4_2 _21649_ (.A(iX[15]),
    .B(iY[15]),
    .C(iX[16]),
    .D(iY[16]),
    .X(_11241_));
 sky130_fd_sc_hd__o21ba_2 _21650_ (.A1(_11017_),
    .A2(_11019_),
    .B1_N(_11015_),
    .X(_11242_));
 sky130_fd_sc_hd__and4_2 _21651_ (.A(iY[15]),
    .B(iX[16]),
    .C(iY[16]),
    .D(iX[17]),
    .X(_11243_));
 sky130_fd_sc_hd__a22oi_2 _21652_ (.A1(iX[16]),
    .A2(iY[16]),
    .B1(iX[17]),
    .B2(iY[15]),
    .Y(_11244_));
 sky130_fd_sc_hd__and4bb_2 _21653_ (.A_N(_11243_),
    .B_N(_11244_),
    .C(iX[15]),
    .D(iY[17]),
    .X(_11246_));
 sky130_fd_sc_hd__o2bb2a_2 _21654_ (.A1_N(iX[15]),
    .A2_N(iY[17]),
    .B1(_11243_),
    .B2(_11244_),
    .X(_11247_));
 sky130_fd_sc_hd__nor2_2 _21655_ (.A(_11246_),
    .B(_11247_),
    .Y(_11248_));
 sky130_fd_sc_hd__xnor2_2 _21656_ (.A(_11242_),
    .B(_11248_),
    .Y(_11249_));
 sky130_fd_sc_hd__o21ai_2 _21657_ (.A1(_11241_),
    .A2(_11101_),
    .B1(_11249_),
    .Y(_11250_));
 sky130_fd_sc_hd__or3_2 _21658_ (.A(_11241_),
    .B(_11101_),
    .C(_11249_),
    .X(_11251_));
 sky130_fd_sc_hd__nand2_2 _21659_ (.A(_11250_),
    .B(_11251_),
    .Y(_11252_));
 sky130_fd_sc_hd__a21oi_2 _21660_ (.A1(_11240_),
    .A2(_11104_),
    .B1(_11252_),
    .Y(_11253_));
 sky130_fd_sc_hd__and3_2 _21661_ (.A(_11240_),
    .B(_11104_),
    .C(_11252_),
    .X(_11254_));
 sky130_fd_sc_hd__nand2_2 _21662_ (.A(iX[12]),
    .B(iY[20]),
    .Y(_11255_));
 sky130_fd_sc_hd__and4_2 _21663_ (.A(iX[13]),
    .B(iX[14]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_11257_));
 sky130_fd_sc_hd__a22oi_2 _21664_ (.A1(iX[14]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[13]),
    .Y(_11258_));
 sky130_fd_sc_hd__nor2_2 _21665_ (.A(_11257_),
    .B(_11258_),
    .Y(_11259_));
 sky130_fd_sc_hd__xnor2_2 _21666_ (.A(_11255_),
    .B(_11259_),
    .Y(_11260_));
 sky130_fd_sc_hd__o21ba_2 _21667_ (.A1(_11084_),
    .A2(_11086_),
    .B1_N(_11083_),
    .X(_11261_));
 sky130_fd_sc_hd__xnor2_2 _21668_ (.A(_11260_),
    .B(_11261_),
    .Y(_11262_));
 sky130_fd_sc_hd__and4_2 _21669_ (.A(iX[10]),
    .B(iX[11]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_11263_));
 sky130_fd_sc_hd__a22oi_2 _21670_ (.A1(iX[11]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[10]),
    .Y(_11264_));
 sky130_fd_sc_hd__nor2_2 _21671_ (.A(_11263_),
    .B(_11264_),
    .Y(_11265_));
 sky130_fd_sc_hd__nand2_2 _21672_ (.A(iX[9]),
    .B(iY[23]),
    .Y(_11266_));
 sky130_fd_sc_hd__xnor2_2 _21673_ (.A(_11265_),
    .B(_11266_),
    .Y(_11268_));
 sky130_fd_sc_hd__and2_2 _21674_ (.A(_11262_),
    .B(_11268_),
    .X(_11269_));
 sky130_fd_sc_hd__nor2_2 _21675_ (.A(_11262_),
    .B(_11268_),
    .Y(_11270_));
 sky130_fd_sc_hd__or2_2 _21676_ (.A(_11269_),
    .B(_11270_),
    .X(_11271_));
 sky130_fd_sc_hd__or3_2 _21677_ (.A(_11253_),
    .B(_11254_),
    .C(_11271_),
    .X(_11272_));
 sky130_fd_sc_hd__o21ai_2 _21678_ (.A1(_11253_),
    .A2(_11254_),
    .B1(_11271_),
    .Y(_11273_));
 sky130_fd_sc_hd__nand3_2 _21679_ (.A(_11239_),
    .B(_11272_),
    .C(_11273_),
    .Y(_11274_));
 sky130_fd_sc_hd__a21o_2 _21680_ (.A1(_11272_),
    .A2(_11273_),
    .B1(_11239_),
    .X(_11275_));
 sky130_fd_sc_hd__nand2_2 _21681_ (.A(_11274_),
    .B(_11275_),
    .Y(_11276_));
 sky130_fd_sc_hd__nor2_2 _21682_ (.A(_11107_),
    .B(_11109_),
    .Y(_11277_));
 sky130_fd_sc_hd__xnor2_2 _21683_ (.A(_11276_),
    .B(_11277_),
    .Y(_11279_));
 sky130_fd_sc_hd__or3_2 _21684_ (.A(_11054_),
    .B(_11058_),
    .C(_11059_),
    .X(_11280_));
 sky130_fd_sc_hd__or2b_2 _21685_ (.A(_11053_),
    .B_N(_11062_),
    .X(_11281_));
 sky130_fd_sc_hd__nand2_2 _21686_ (.A(iY[11]),
    .B(iX[21]),
    .Y(_11282_));
 sky130_fd_sc_hd__and4_2 _21687_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[22]),
    .D(iX[23]),
    .X(_11283_));
 sky130_fd_sc_hd__a22oi_2 _21688_ (.A1(iY[10]),
    .A2(iX[22]),
    .B1(iX[23]),
    .B2(iY[9]),
    .Y(_11284_));
 sky130_fd_sc_hd__nor2_2 _21689_ (.A(_11283_),
    .B(_11284_),
    .Y(_11285_));
 sky130_fd_sc_hd__xnor2_2 _21690_ (.A(_11282_),
    .B(_11285_),
    .Y(_11286_));
 sky130_fd_sc_hd__o21ba_2 _21691_ (.A1(_11022_),
    .A2(_11024_),
    .B1_N(_11021_),
    .X(_11287_));
 sky130_fd_sc_hd__xnor2_2 _21692_ (.A(_11286_),
    .B(_11287_),
    .Y(_11288_));
 sky130_fd_sc_hd__nand2_2 _21693_ (.A(iY[14]),
    .B(iX[18]),
    .Y(_11290_));
 sky130_fd_sc_hd__and4_2 _21694_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[19]),
    .D(iX[20]),
    .X(_11291_));
 sky130_fd_sc_hd__a22oi_2 _21695_ (.A1(iY[13]),
    .A2(iX[19]),
    .B1(iX[20]),
    .B2(iY[12]),
    .Y(_11292_));
 sky130_fd_sc_hd__nor2_2 _21696_ (.A(_11291_),
    .B(_11292_),
    .Y(_11293_));
 sky130_fd_sc_hd__xnor2_2 _21697_ (.A(_11290_),
    .B(_11293_),
    .Y(_11294_));
 sky130_fd_sc_hd__and2_2 _21698_ (.A(_11288_),
    .B(_11294_),
    .X(_11295_));
 sky130_fd_sc_hd__nor2_2 _21699_ (.A(_11288_),
    .B(_11294_),
    .Y(_11296_));
 sky130_fd_sc_hd__or2_2 _21700_ (.A(_11295_),
    .B(_11296_),
    .X(_11297_));
 sky130_fd_sc_hd__a21o_2 _21701_ (.A1(_11280_),
    .A2(_11281_),
    .B1(_11297_),
    .X(_11298_));
 sky130_fd_sc_hd__nand3_2 _21702_ (.A(_11280_),
    .B(_11281_),
    .C(_11297_),
    .Y(_11299_));
 sky130_fd_sc_hd__and2b_2 _21703_ (.A_N(_11026_),
    .B(_11025_),
    .X(_11301_));
 sky130_fd_sc_hd__a21o_2 _21704_ (.A1(_11020_),
    .A2(_11028_),
    .B1(_11301_),
    .X(_11302_));
 sky130_fd_sc_hd__a21o_2 _21705_ (.A1(_11298_),
    .A2(_11299_),
    .B1(_11302_),
    .X(_11303_));
 sky130_fd_sc_hd__nand3_2 _21706_ (.A(_11298_),
    .B(_11299_),
    .C(_11302_),
    .Y(_11304_));
 sky130_fd_sc_hd__and2_2 _21707_ (.A(_11303_),
    .B(_11304_),
    .X(_11305_));
 sky130_fd_sc_hd__and4_2 _21708_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[25]),
    .D(iX[26]),
    .X(_11306_));
 sky130_fd_sc_hd__a22oi_2 _21709_ (.A1(iY[7]),
    .A2(iX[25]),
    .B1(iX[26]),
    .B2(iY[6]),
    .Y(_11307_));
 sky130_fd_sc_hd__and4bb_2 _21710_ (.A_N(_11306_),
    .B_N(_11307_),
    .C(iY[8]),
    .D(iX[24]),
    .X(_11308_));
 sky130_fd_sc_hd__o2bb2a_2 _21711_ (.A1_N(iY[8]),
    .A2_N(iX[24]),
    .B1(_11306_),
    .B2(_11307_),
    .X(_11309_));
 sky130_fd_sc_hd__nor2_2 _21712_ (.A(_11308_),
    .B(_11309_),
    .Y(_11310_));
 sky130_fd_sc_hd__o21ai_2 _21713_ (.A1(_11043_),
    .A2(_11047_),
    .B1(_11310_),
    .Y(_11311_));
 sky130_fd_sc_hd__or3_2 _21714_ (.A(_11043_),
    .B(_11047_),
    .C(_11310_),
    .X(_11312_));
 sky130_fd_sc_hd__and2_2 _21715_ (.A(_11311_),
    .B(_11312_),
    .X(_11313_));
 sky130_fd_sc_hd__or3_2 _21716_ (.A(_11055_),
    .B(_11059_),
    .C(_11313_),
    .X(_11314_));
 sky130_fd_sc_hd__o21ai_2 _21717_ (.A1(_11055_),
    .A2(_11059_),
    .B1(_11313_),
    .Y(_11315_));
 sky130_fd_sc_hd__nand2_2 _21718_ (.A(_11314_),
    .B(_11315_),
    .Y(_11316_));
 sky130_fd_sc_hd__nand2_2 _21719_ (.A(_11040_),
    .B(_11041_),
    .Y(_11317_));
 sky130_fd_sc_hd__or3_2 _21720_ (.A(_11042_),
    .B(_11046_),
    .C(_11047_),
    .X(_11318_));
 sky130_fd_sc_hd__and4_2 _21721_ (.A(iY[3]),
    .B(iY[4]),
    .C(iX[28]),
    .D(iX[29]),
    .X(_11319_));
 sky130_fd_sc_hd__a22oi_2 _21722_ (.A1(iY[4]),
    .A2(iX[28]),
    .B1(iX[29]),
    .B2(iY[3]),
    .Y(_11320_));
 sky130_fd_sc_hd__nor2_2 _21723_ (.A(_11319_),
    .B(_11320_),
    .Y(_11322_));
 sky130_fd_sc_hd__nand2_2 _21724_ (.A(iY[5]),
    .B(iX[27]),
    .Y(_11323_));
 sky130_fd_sc_hd__xnor2_2 _21725_ (.A(_11322_),
    .B(_11323_),
    .Y(_11324_));
 sky130_fd_sc_hd__and4_2 _21726_ (.A(iY[1]),
    .B(iY[2]),
    .C(iX[30]),
    .D(iX[31]),
    .X(_11325_));
 sky130_fd_sc_hd__a22oi_2 _21727_ (.A1(iY[2]),
    .A2(iX[30]),
    .B1(iX[31]),
    .B2(iY[1]),
    .Y(_11326_));
 sky130_fd_sc_hd__or2_2 _21728_ (.A(_11325_),
    .B(_11326_),
    .X(_11327_));
 sky130_fd_sc_hd__a31o_2 _21729_ (.A1(iY[2]),
    .A2(iX[29]),
    .A3(_11037_),
    .B1(_11036_),
    .X(_11328_));
 sky130_fd_sc_hd__xnor2_2 _21730_ (.A(_11327_),
    .B(_11328_),
    .Y(_11329_));
 sky130_fd_sc_hd__xnor2_2 _21731_ (.A(_11324_),
    .B(_11329_),
    .Y(_11330_));
 sky130_fd_sc_hd__a21oi_2 _21732_ (.A1(_11317_),
    .A2(_11318_),
    .B1(_11330_),
    .Y(_11331_));
 sky130_fd_sc_hd__and3_2 _21733_ (.A(_11317_),
    .B(_11318_),
    .C(_11330_),
    .X(_11333_));
 sky130_fd_sc_hd__or2_2 _21734_ (.A(_11331_),
    .B(_11333_),
    .X(_11334_));
 sky130_fd_sc_hd__nor2_2 _21735_ (.A(_11316_),
    .B(_11334_),
    .Y(_11335_));
 sky130_fd_sc_hd__and2_2 _21736_ (.A(_11316_),
    .B(_11334_),
    .X(_11336_));
 sky130_fd_sc_hd__or2_2 _21737_ (.A(_11335_),
    .B(_11336_),
    .X(_11337_));
 sky130_fd_sc_hd__and2_2 _21738_ (.A(_11051_),
    .B(_11064_),
    .X(_11338_));
 sky130_fd_sc_hd__xor2_2 _21739_ (.A(_11337_),
    .B(_11338_),
    .X(_11339_));
 sky130_fd_sc_hd__nand2_2 _21740_ (.A(_11305_),
    .B(_11339_),
    .Y(_11340_));
 sky130_fd_sc_hd__or2_2 _21741_ (.A(_11305_),
    .B(_11339_),
    .X(_11341_));
 sky130_fd_sc_hd__o211a_2 _21742_ (.A1(_11067_),
    .A2(_11072_),
    .B1(_11340_),
    .C1(_11341_),
    .X(_11342_));
 sky130_fd_sc_hd__nand2_2 _21743_ (.A(_11340_),
    .B(_11341_),
    .Y(_11344_));
 sky130_fd_sc_hd__or3b_2 _21744_ (.A(_11067_),
    .B(_11072_),
    .C_N(_11344_),
    .X(_11345_));
 sky130_fd_sc_hd__or2b_2 _21745_ (.A(_11342_),
    .B_N(_11345_),
    .X(_11346_));
 sky130_fd_sc_hd__xor2_2 _21746_ (.A(_11279_),
    .B(_11346_),
    .X(_11347_));
 sky130_fd_sc_hd__o21ai_2 _21747_ (.A1(_11074_),
    .A2(_11116_),
    .B1(_11347_),
    .Y(_11348_));
 sky130_fd_sc_hd__or3_2 _21748_ (.A(_11074_),
    .B(_11116_),
    .C(_11347_),
    .X(_11349_));
 sky130_fd_sc_hd__and2_2 _21749_ (.A(_11348_),
    .B(_11349_),
    .X(_11350_));
 sky130_fd_sc_hd__nand2_2 _21750_ (.A(_11238_),
    .B(_11350_),
    .Y(_11351_));
 sky130_fd_sc_hd__or2_2 _21751_ (.A(_11238_),
    .B(_11350_),
    .X(_11352_));
 sky130_fd_sc_hd__nand2_2 _21752_ (.A(_11351_),
    .B(_11352_),
    .Y(_11353_));
 sky130_fd_sc_hd__a21o_2 _21753_ (.A1(_11118_),
    .A2(_11171_),
    .B1(_11353_),
    .X(_11355_));
 sky130_fd_sc_hd__nand3_2 _21754_ (.A(_11118_),
    .B(_11171_),
    .C(_11353_),
    .Y(_11356_));
 sky130_fd_sc_hd__nand2_2 _21755_ (.A(_11355_),
    .B(_11356_),
    .Y(_11357_));
 sky130_fd_sc_hd__xor2_2 _21756_ (.A(_11192_),
    .B(_11357_),
    .X(_11358_));
 sky130_fd_sc_hd__and2_2 _21757_ (.A(_11173_),
    .B(_11175_),
    .X(_11359_));
 sky130_fd_sc_hd__or2_2 _21758_ (.A(_11358_),
    .B(_11359_),
    .X(_11360_));
 sky130_fd_sc_hd__nand2_2 _21759_ (.A(_11358_),
    .B(_11359_),
    .Y(_11361_));
 sky130_fd_sc_hd__nand2_2 _21760_ (.A(_11360_),
    .B(_11361_),
    .Y(_11362_));
 sky130_fd_sc_hd__xnor2_2 _21761_ (.A(_11191_),
    .B(_11362_),
    .Y(_11363_));
 sky130_fd_sc_hd__o21a_2 _21762_ (.A1(_11189_),
    .A2(_11181_),
    .B1(_11363_),
    .X(_11364_));
 sky130_fd_sc_hd__nor3_2 _21763_ (.A(_11189_),
    .B(_11181_),
    .C(_11363_),
    .Y(_11366_));
 sky130_fd_sc_hd__or2_2 _21764_ (.A(_11364_),
    .B(_11366_),
    .X(_11367_));
 sky130_fd_sc_hd__a21oi_2 _21765_ (.A1(_11188_),
    .A2(_11185_),
    .B1(_11367_),
    .Y(_11368_));
 sky130_fd_sc_hd__and3_2 _21766_ (.A(_11188_),
    .B(_11185_),
    .C(_11367_),
    .X(_11369_));
 sky130_fd_sc_hd__or2_2 _21767_ (.A(_11368_),
    .B(_11369_),
    .X(_11370_));
 sky130_fd_sc_hd__nand2_2 _21768_ (.A(iX[0]),
    .B(iX[32]),
    .Y(_11371_));
 sky130_fd_sc_hd__or2_2 _21769_ (.A(iX[0]),
    .B(iX[32]),
    .X(_11372_));
 sky130_fd_sc_hd__and2_2 _21770_ (.A(_11371_),
    .B(_11372_),
    .X(_11373_));
 sky130_fd_sc_hd__buf_6 _21771_ (.A(_11373_),
    .X(_11374_));
 sky130_fd_sc_hd__nand2_2 _21772_ (.A(iY[0]),
    .B(iY[32]),
    .Y(_11375_));
 sky130_fd_sc_hd__or2_2 _21773_ (.A(iY[0]),
    .B(iY[32]),
    .X(_11377_));
 sky130_fd_sc_hd__and2_2 _21774_ (.A(_11375_),
    .B(_11377_),
    .X(_11378_));
 sky130_fd_sc_hd__buf_1 _21775_ (.A(_11378_),
    .X(_11379_));
 sky130_fd_sc_hd__buf_4 _21776_ (.A(_11379_),
    .X(_11380_));
 sky130_fd_sc_hd__buf_2 _21777_ (.A(_11380_),
    .X(_11381_));
 sky130_fd_sc_hd__nand2_2 _21778_ (.A(_11374_),
    .B(_11381_),
    .Y(_11382_));
 sky130_fd_sc_hd__nand2_2 _21779_ (.A(iX[32]),
    .B(iY[32]),
    .Y(_11383_));
 sky130_fd_sc_hd__xor2_2 _21780_ (.A(_11382_),
    .B(_11383_),
    .X(_11384_));
 sky130_fd_sc_hd__xnor2_2 _21781_ (.A(_10801_),
    .B(_11384_),
    .Y(_11385_));
 sky130_fd_sc_hd__and2b_2 _21782_ (.A_N(_11370_),
    .B(_11385_),
    .X(_11386_));
 sky130_fd_sc_hd__or2b_2 _21783_ (.A(_11362_),
    .B_N(_11191_),
    .X(_11388_));
 sky130_fd_sc_hd__or2b_2 _21784_ (.A(_11357_),
    .B_N(_11192_),
    .X(_11389_));
 sky130_fd_sc_hd__or2b_2 _21785_ (.A(_11236_),
    .B_N(_11237_),
    .X(_11390_));
 sky130_fd_sc_hd__nor2_2 _21786_ (.A(_11279_),
    .B(_11346_),
    .Y(_11391_));
 sky130_fd_sc_hd__or2_2 _21787_ (.A(_11337_),
    .B(_11338_),
    .X(_11392_));
 sky130_fd_sc_hd__nand2_2 _21788_ (.A(iY[1]),
    .B(iX[30]),
    .Y(_11393_));
 sky130_fd_sc_hd__and3_2 _21789_ (.A(iY[2]),
    .B(iX[31]),
    .C(_11393_),
    .X(_11394_));
 sky130_fd_sc_hd__and2_2 _21790_ (.A(iY[4]),
    .B(iX[30]),
    .X(_11395_));
 sky130_fd_sc_hd__nand3_2 _21791_ (.A(iY[3]),
    .B(iX[29]),
    .C(_11395_),
    .Y(_11396_));
 sky130_fd_sc_hd__a22o_2 _21792_ (.A1(iY[4]),
    .A2(iX[29]),
    .B1(iX[30]),
    .B2(iY[3]),
    .X(_11397_));
 sky130_fd_sc_hd__and2_2 _21793_ (.A(iY[5]),
    .B(iX[28]),
    .X(_11399_));
 sky130_fd_sc_hd__a21oi_2 _21794_ (.A1(_11396_),
    .A2(_11397_),
    .B1(_11399_),
    .Y(_11400_));
 sky130_fd_sc_hd__and3_2 _21795_ (.A(_11396_),
    .B(_11397_),
    .C(_11399_),
    .X(_11401_));
 sky130_fd_sc_hd__nor2_2 _21796_ (.A(_11400_),
    .B(_11401_),
    .Y(_11402_));
 sky130_fd_sc_hd__xnor2_2 _21797_ (.A(_11394_),
    .B(_11402_),
    .Y(_11403_));
 sky130_fd_sc_hd__or2b_2 _21798_ (.A(_11327_),
    .B_N(_11328_),
    .X(_11404_));
 sky130_fd_sc_hd__a21bo_2 _21799_ (.A1(_11324_),
    .A2(_11329_),
    .B1_N(_11404_),
    .X(_11405_));
 sky130_fd_sc_hd__xor2_2 _21800_ (.A(_11403_),
    .B(_11405_),
    .X(_11406_));
 sky130_fd_sc_hd__o21ba_2 _21801_ (.A1(_11320_),
    .A2(_11323_),
    .B1_N(_11319_),
    .X(_11407_));
 sky130_fd_sc_hd__and4_2 _21802_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[26]),
    .D(iX[27]),
    .X(_11408_));
 sky130_fd_sc_hd__a22oi_2 _21803_ (.A1(iY[7]),
    .A2(iX[26]),
    .B1(iX[27]),
    .B2(iY[6]),
    .Y(_11410_));
 sky130_fd_sc_hd__nor2_2 _21804_ (.A(_11408_),
    .B(_11410_),
    .Y(_11411_));
 sky130_fd_sc_hd__nand2_2 _21805_ (.A(iY[8]),
    .B(iX[25]),
    .Y(_11412_));
 sky130_fd_sc_hd__xnor2_2 _21806_ (.A(_11411_),
    .B(_11412_),
    .Y(_11413_));
 sky130_fd_sc_hd__xnor2_2 _21807_ (.A(_11407_),
    .B(_11413_),
    .Y(_11414_));
 sky130_fd_sc_hd__o21ai_2 _21808_ (.A1(_11306_),
    .A2(_11308_),
    .B1(_11414_),
    .Y(_11415_));
 sky130_fd_sc_hd__or3_2 _21809_ (.A(_11306_),
    .B(_11308_),
    .C(_11414_),
    .X(_11416_));
 sky130_fd_sc_hd__nand2_2 _21810_ (.A(_11415_),
    .B(_11416_),
    .Y(_11417_));
 sky130_fd_sc_hd__nor2_2 _21811_ (.A(_11406_),
    .B(_11417_),
    .Y(_11418_));
 sky130_fd_sc_hd__and2_2 _21812_ (.A(_11406_),
    .B(_11417_),
    .X(_11419_));
 sky130_fd_sc_hd__nor2_2 _21813_ (.A(_11418_),
    .B(_11419_),
    .Y(_11421_));
 sky130_fd_sc_hd__o21a_2 _21814_ (.A1(_11331_),
    .A2(_11335_),
    .B1(_11421_),
    .X(_11422_));
 sky130_fd_sc_hd__nor3_2 _21815_ (.A(_11331_),
    .B(_11335_),
    .C(_11421_),
    .Y(_11423_));
 sky130_fd_sc_hd__nor2_2 _21816_ (.A(_11422_),
    .B(_11423_),
    .Y(_11424_));
 sky130_fd_sc_hd__and2b_2 _21817_ (.A_N(_11287_),
    .B(_11286_),
    .X(_11425_));
 sky130_fd_sc_hd__and4_2 _21818_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[20]),
    .D(iX[21]),
    .X(_11426_));
 sky130_fd_sc_hd__a22oi_2 _21819_ (.A1(iY[13]),
    .A2(iX[20]),
    .B1(iX[21]),
    .B2(iY[12]),
    .Y(_11427_));
 sky130_fd_sc_hd__nor2_2 _21820_ (.A(_11426_),
    .B(_11427_),
    .Y(_11428_));
 sky130_fd_sc_hd__nand2_2 _21821_ (.A(iY[14]),
    .B(iX[19]),
    .Y(_11429_));
 sky130_fd_sc_hd__xnor2_2 _21822_ (.A(_11428_),
    .B(_11429_),
    .Y(_11430_));
 sky130_fd_sc_hd__and4_2 _21823_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[23]),
    .D(iX[24]),
    .X(_11432_));
 sky130_fd_sc_hd__a22oi_2 _21824_ (.A1(iY[10]),
    .A2(iX[23]),
    .B1(iX[24]),
    .B2(iY[9]),
    .Y(_11433_));
 sky130_fd_sc_hd__nor2_2 _21825_ (.A(_11432_),
    .B(_11433_),
    .Y(_11434_));
 sky130_fd_sc_hd__nand2_2 _21826_ (.A(iY[11]),
    .B(iX[22]),
    .Y(_11435_));
 sky130_fd_sc_hd__xnor2_2 _21827_ (.A(_11434_),
    .B(_11435_),
    .Y(_11436_));
 sky130_fd_sc_hd__o21ba_2 _21828_ (.A1(_11282_),
    .A2(_11284_),
    .B1_N(_11283_),
    .X(_11437_));
 sky130_fd_sc_hd__xnor2_2 _21829_ (.A(_11436_),
    .B(_11437_),
    .Y(_11438_));
 sky130_fd_sc_hd__xnor2_2 _21830_ (.A(_11430_),
    .B(_11438_),
    .Y(_11439_));
 sky130_fd_sc_hd__a21o_2 _21831_ (.A1(_11311_),
    .A2(_11315_),
    .B1(_11439_),
    .X(_11440_));
 sky130_fd_sc_hd__nand3_2 _21832_ (.A(_11311_),
    .B(_11315_),
    .C(_11439_),
    .Y(_11441_));
 sky130_fd_sc_hd__o211ai_2 _21833_ (.A1(_11425_),
    .A2(_11295_),
    .B1(_11440_),
    .C1(_11441_),
    .Y(_11443_));
 sky130_fd_sc_hd__a211o_2 _21834_ (.A1(_11440_),
    .A2(_11441_),
    .B1(_11425_),
    .C1(_11295_),
    .X(_11444_));
 sky130_fd_sc_hd__and2_2 _21835_ (.A(_11443_),
    .B(_11444_),
    .X(_11445_));
 sky130_fd_sc_hd__xnor2_2 _21836_ (.A(_11424_),
    .B(_11445_),
    .Y(_11446_));
 sky130_fd_sc_hd__a21oi_2 _21837_ (.A1(_11392_),
    .A2(_11340_),
    .B1(_11446_),
    .Y(_11447_));
 sky130_fd_sc_hd__and3_2 _21838_ (.A(_11392_),
    .B(_11340_),
    .C(_11446_),
    .X(_11448_));
 sky130_fd_sc_hd__or2_2 _21839_ (.A(_11447_),
    .B(_11448_),
    .X(_11449_));
 sky130_fd_sc_hd__or2b_2 _21840_ (.A(_11253_),
    .B_N(_11272_),
    .X(_11450_));
 sky130_fd_sc_hd__and4_2 _21841_ (.A(iX[11]),
    .B(iX[12]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_11451_));
 sky130_fd_sc_hd__a22oi_2 _21842_ (.A1(iX[12]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[11]),
    .Y(_11452_));
 sky130_fd_sc_hd__nor2_2 _21843_ (.A(_11451_),
    .B(_11452_),
    .Y(_11454_));
 sky130_fd_sc_hd__nand2_2 _21844_ (.A(iX[10]),
    .B(iY[23]),
    .Y(_11455_));
 sky130_fd_sc_hd__xnor2_2 _21845_ (.A(_11454_),
    .B(_11455_),
    .Y(_11456_));
 sky130_fd_sc_hd__and4_2 _21846_ (.A(iX[14]),
    .B(iX[15]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_11457_));
 sky130_fd_sc_hd__a22oi_2 _21847_ (.A1(iX[15]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[14]),
    .Y(_11458_));
 sky130_fd_sc_hd__nor2_2 _21848_ (.A(_11457_),
    .B(_11458_),
    .Y(_11459_));
 sky130_fd_sc_hd__nand2_2 _21849_ (.A(iX[13]),
    .B(iY[20]),
    .Y(_11460_));
 sky130_fd_sc_hd__xnor2_2 _21850_ (.A(_11459_),
    .B(_11460_),
    .Y(_11461_));
 sky130_fd_sc_hd__o21ba_2 _21851_ (.A1(_11255_),
    .A2(_11258_),
    .B1_N(_11257_),
    .X(_11462_));
 sky130_fd_sc_hd__xnor2_2 _21852_ (.A(_11461_),
    .B(_11462_),
    .Y(_11463_));
 sky130_fd_sc_hd__and2_2 _21853_ (.A(_11456_),
    .B(_11463_),
    .X(_11465_));
 sky130_fd_sc_hd__nor2_2 _21854_ (.A(_11456_),
    .B(_11463_),
    .Y(_11466_));
 sky130_fd_sc_hd__or2_2 _21855_ (.A(_11465_),
    .B(_11466_),
    .X(_11467_));
 sky130_fd_sc_hd__or3_2 _21856_ (.A(_11242_),
    .B(_11246_),
    .C(_11247_),
    .X(_11468_));
 sky130_fd_sc_hd__o21ba_2 _21857_ (.A1(_11290_),
    .A2(_11292_),
    .B1_N(_11291_),
    .X(_11469_));
 sky130_fd_sc_hd__and4_2 _21858_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[17]),
    .D(iX[18]),
    .X(_11470_));
 sky130_fd_sc_hd__a22oi_2 _21859_ (.A1(iY[16]),
    .A2(iX[17]),
    .B1(iX[18]),
    .B2(iY[15]),
    .Y(_11471_));
 sky130_fd_sc_hd__and4bb_2 _21860_ (.A_N(_11470_),
    .B_N(_11471_),
    .C(iX[16]),
    .D(iY[17]),
    .X(_11472_));
 sky130_fd_sc_hd__o2bb2a_2 _21861_ (.A1_N(iX[16]),
    .A2_N(iY[17]),
    .B1(_11470_),
    .B2(_11471_),
    .X(_11473_));
 sky130_fd_sc_hd__nor2_2 _21862_ (.A(_11472_),
    .B(_11473_),
    .Y(_11474_));
 sky130_fd_sc_hd__xnor2_2 _21863_ (.A(_11469_),
    .B(_11474_),
    .Y(_11476_));
 sky130_fd_sc_hd__o21ai_2 _21864_ (.A1(_11243_),
    .A2(_11246_),
    .B1(_11476_),
    .Y(_11477_));
 sky130_fd_sc_hd__or3_2 _21865_ (.A(_11243_),
    .B(_11246_),
    .C(_11476_),
    .X(_11478_));
 sky130_fd_sc_hd__nand2_2 _21866_ (.A(_11477_),
    .B(_11478_),
    .Y(_11479_));
 sky130_fd_sc_hd__a21oi_2 _21867_ (.A1(_11468_),
    .A2(_11250_),
    .B1(_11479_),
    .Y(_11480_));
 sky130_fd_sc_hd__and3_2 _21868_ (.A(_11468_),
    .B(_11250_),
    .C(_11479_),
    .X(_11481_));
 sky130_fd_sc_hd__or3_2 _21869_ (.A(_11467_),
    .B(_11480_),
    .C(_11481_),
    .X(_11482_));
 sky130_fd_sc_hd__o21ai_2 _21870_ (.A1(_11480_),
    .A2(_11481_),
    .B1(_11467_),
    .Y(_11483_));
 sky130_fd_sc_hd__nand2_2 _21871_ (.A(_11482_),
    .B(_11483_),
    .Y(_11484_));
 sky130_fd_sc_hd__a21oi_2 _21872_ (.A1(_11298_),
    .A2(_11304_),
    .B1(_11484_),
    .Y(_11485_));
 sky130_fd_sc_hd__and3_2 _21873_ (.A(_11298_),
    .B(_11304_),
    .C(_11484_),
    .X(_11487_));
 sky130_fd_sc_hd__nor2_2 _21874_ (.A(_11485_),
    .B(_11487_),
    .Y(_11488_));
 sky130_fd_sc_hd__xnor2_2 _21875_ (.A(_11450_),
    .B(_11488_),
    .Y(_11489_));
 sky130_fd_sc_hd__nor2_2 _21876_ (.A(_11449_),
    .B(_11489_),
    .Y(_11490_));
 sky130_fd_sc_hd__and2_2 _21877_ (.A(_11449_),
    .B(_11489_),
    .X(_11491_));
 sky130_fd_sc_hd__nor2_2 _21878_ (.A(_11490_),
    .B(_11491_),
    .Y(_11492_));
 sky130_fd_sc_hd__o21a_2 _21879_ (.A1(_11342_),
    .A2(_11391_),
    .B1(_11492_),
    .X(_11493_));
 sky130_fd_sc_hd__nor3_2 _21880_ (.A(_11342_),
    .B(_11391_),
    .C(_11492_),
    .Y(_11494_));
 sky130_fd_sc_hd__nor2_2 _21881_ (.A(_11493_),
    .B(_11494_),
    .Y(_11495_));
 sky130_fd_sc_hd__a21boi_2 _21882_ (.A1(_11213_),
    .A2(_11229_),
    .B1_N(_11211_),
    .Y(_11496_));
 sky130_fd_sc_hd__o21a_2 _21883_ (.A1(_11276_),
    .A2(_11277_),
    .B1(_11274_),
    .X(_11498_));
 sky130_fd_sc_hd__or2b_2 _21884_ (.A(_11220_),
    .B_N(_11219_),
    .X(_11499_));
 sky130_fd_sc_hd__and4_2 _21885_ (.A(iX[5]),
    .B(iX[6]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_11500_));
 sky130_fd_sc_hd__a22oi_2 _21886_ (.A1(iX[6]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[5]),
    .Y(_11501_));
 sky130_fd_sc_hd__nor2_2 _21887_ (.A(_11500_),
    .B(_11501_),
    .Y(_11502_));
 sky130_fd_sc_hd__nand2_2 _21888_ (.A(iX[4]),
    .B(iY[29]),
    .Y(_11503_));
 sky130_fd_sc_hd__xnor2_2 _21889_ (.A(_11502_),
    .B(_11503_),
    .Y(_11504_));
 sky130_fd_sc_hd__o21ba_2 _21890_ (.A1(_11215_),
    .A2(_11217_),
    .B1_N(_11216_),
    .X(_11505_));
 sky130_fd_sc_hd__xnor2_2 _21891_ (.A(_11504_),
    .B(_11505_),
    .Y(_11506_));
 sky130_fd_sc_hd__nand3_2 _21892_ (.A(iX[3]),
    .B(iY[30]),
    .C(_11506_),
    .Y(_11507_));
 sky130_fd_sc_hd__a21o_2 _21893_ (.A1(iX[3]),
    .A2(iY[30]),
    .B1(_11506_),
    .X(_11509_));
 sky130_fd_sc_hd__nand2_2 _21894_ (.A(_11507_),
    .B(_11509_),
    .Y(_11510_));
 sky130_fd_sc_hd__a21oi_2 _21895_ (.A1(_11499_),
    .A2(_11222_),
    .B1(_11510_),
    .Y(_11511_));
 sky130_fd_sc_hd__and3_2 _21896_ (.A(_11499_),
    .B(_11222_),
    .C(_11510_),
    .X(_11512_));
 sky130_fd_sc_hd__nor2_2 _21897_ (.A(_11511_),
    .B(_11512_),
    .Y(_11513_));
 sky130_fd_sc_hd__nand2_2 _21898_ (.A(iX[2]),
    .B(iY[31]),
    .Y(_11514_));
 sky130_fd_sc_hd__xnor2_2 _21899_ (.A(_11513_),
    .B(_11514_),
    .Y(_11515_));
 sky130_fd_sc_hd__and2b_2 _21900_ (.A_N(_11209_),
    .B(_11195_),
    .X(_11516_));
 sky130_fd_sc_hd__or2b_2 _21901_ (.A(_11198_),
    .B_N(_11204_),
    .X(_11517_));
 sky130_fd_sc_hd__or2b_2 _21902_ (.A(_11197_),
    .B_N(_11205_),
    .X(_11518_));
 sky130_fd_sc_hd__nand2_2 _21903_ (.A(_11517_),
    .B(_11518_),
    .Y(_11520_));
 sky130_fd_sc_hd__and2b_2 _21904_ (.A_N(_11261_),
    .B(_11260_),
    .X(_11521_));
 sky130_fd_sc_hd__o21ba_2 _21905_ (.A1(_11199_),
    .A2(_11202_),
    .B1_N(_11200_),
    .X(_11522_));
 sky130_fd_sc_hd__o21ba_2 _21906_ (.A1(_11264_),
    .A2(_11266_),
    .B1_N(_11263_),
    .X(_11523_));
 sky130_fd_sc_hd__and4_2 _21907_ (.A(iX[8]),
    .B(iX[9]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_11524_));
 sky130_fd_sc_hd__a22oi_2 _21908_ (.A1(iX[9]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[8]),
    .Y(_11525_));
 sky130_fd_sc_hd__nor2_2 _21909_ (.A(_11524_),
    .B(_11525_),
    .Y(_11526_));
 sky130_fd_sc_hd__nand2_2 _21910_ (.A(iX[7]),
    .B(iY[26]),
    .Y(_11527_));
 sky130_fd_sc_hd__xnor2_2 _21911_ (.A(_11526_),
    .B(_11527_),
    .Y(_11528_));
 sky130_fd_sc_hd__xnor2_2 _21912_ (.A(_11523_),
    .B(_11528_),
    .Y(_11529_));
 sky130_fd_sc_hd__xnor2_2 _21913_ (.A(_11522_),
    .B(_11529_),
    .Y(_11530_));
 sky130_fd_sc_hd__o21a_2 _21914_ (.A1(_11521_),
    .A2(_11269_),
    .B1(_11530_),
    .X(_11531_));
 sky130_fd_sc_hd__nor3_2 _21915_ (.A(_11521_),
    .B(_11269_),
    .C(_11530_),
    .Y(_11532_));
 sky130_fd_sc_hd__or2_2 _21916_ (.A(_11531_),
    .B(_11532_),
    .X(_11533_));
 sky130_fd_sc_hd__xnor2_2 _21917_ (.A(_11520_),
    .B(_11533_),
    .Y(_11534_));
 sky130_fd_sc_hd__o21a_2 _21918_ (.A1(_11207_),
    .A2(_11516_),
    .B1(_11534_),
    .X(_11535_));
 sky130_fd_sc_hd__inv_2 _21919_ (.A(_11535_),
    .Y(_11536_));
 sky130_fd_sc_hd__or3_2 _21920_ (.A(_11207_),
    .B(_11516_),
    .C(_11534_),
    .X(_11537_));
 sky130_fd_sc_hd__and3_2 _21921_ (.A(_11515_),
    .B(_11536_),
    .C(_11537_),
    .X(_11538_));
 sky130_fd_sc_hd__a21oi_2 _21922_ (.A1(_11536_),
    .A2(_11537_),
    .B1(_11515_),
    .Y(_11539_));
 sky130_fd_sc_hd__or2_2 _21923_ (.A(_11538_),
    .B(_11539_),
    .X(_11541_));
 sky130_fd_sc_hd__xor2_2 _21924_ (.A(_11498_),
    .B(_11541_),
    .X(_11542_));
 sky130_fd_sc_hd__xnor2_2 _21925_ (.A(_11496_),
    .B(_11542_),
    .Y(_11543_));
 sky130_fd_sc_hd__xnor2_2 _21926_ (.A(_11495_),
    .B(_11543_),
    .Y(_11544_));
 sky130_fd_sc_hd__a21oi_2 _21927_ (.A1(_11348_),
    .A2(_11351_),
    .B1(_11544_),
    .Y(_11545_));
 sky130_fd_sc_hd__and3_2 _21928_ (.A(_11348_),
    .B(_11351_),
    .C(_11544_),
    .X(_11546_));
 sky130_fd_sc_hd__or2_2 _21929_ (.A(_11545_),
    .B(_11546_),
    .X(_11547_));
 sky130_fd_sc_hd__a21oi_2 _21930_ (.A1(_11233_),
    .A2(_11390_),
    .B1(_11547_),
    .Y(_11548_));
 sky130_fd_sc_hd__and3_2 _21931_ (.A(_11233_),
    .B(_11390_),
    .C(_11547_),
    .X(_11549_));
 sky130_fd_sc_hd__or2_2 _21932_ (.A(_11548_),
    .B(_11549_),
    .X(_11550_));
 sky130_fd_sc_hd__a21oi_2 _21933_ (.A1(_11355_),
    .A2(_11389_),
    .B1(_11550_),
    .Y(_11552_));
 sky130_fd_sc_hd__and3_2 _21934_ (.A(_11355_),
    .B(_11389_),
    .C(_11550_),
    .X(_11553_));
 sky130_fd_sc_hd__or2_2 _21935_ (.A(_11552_),
    .B(_11553_),
    .X(_11554_));
 sky130_fd_sc_hd__o21ba_2 _21936_ (.A1(_11214_),
    .A2(_11227_),
    .B1_N(_11226_),
    .X(_11555_));
 sky130_fd_sc_hd__xnor2_2 _21937_ (.A(_11554_),
    .B(_11555_),
    .Y(_11556_));
 sky130_fd_sc_hd__a21oi_2 _21938_ (.A1(_11360_),
    .A2(_11388_),
    .B1(_11556_),
    .Y(_11557_));
 sky130_fd_sc_hd__and3_2 _21939_ (.A(_11360_),
    .B(_11388_),
    .C(_11556_),
    .X(_11558_));
 sky130_fd_sc_hd__or2_2 _21940_ (.A(_11557_),
    .B(_11558_),
    .X(_11559_));
 sky130_fd_sc_hd__o21bai_2 _21941_ (.A1(_11364_),
    .A2(_11368_),
    .B1_N(_11559_),
    .Y(_11560_));
 sky130_fd_sc_hd__or3b_2 _21942_ (.A(_11364_),
    .B(_11368_),
    .C_N(_11559_),
    .X(_11561_));
 sky130_fd_sc_hd__o21a_2 _21943_ (.A1(oO[0]),
    .A2(_11384_),
    .B1(_11382_),
    .X(_11563_));
 sky130_fd_sc_hd__nand2_2 _21944_ (.A(_11375_),
    .B(_11377_),
    .Y(_11564_));
 sky130_fd_sc_hd__buf_1 _21945_ (.A(_11564_),
    .X(_11565_));
 sky130_fd_sc_hd__buf_1 _21946_ (.A(_11565_),
    .X(_11566_));
 sky130_fd_sc_hd__buf_1 _21947_ (.A(_11566_),
    .X(_11567_));
 sky130_fd_sc_hd__xor2_4 _21948_ (.A(iX[1]),
    .B(iX[33]),
    .X(_11568_));
 sky130_fd_sc_hd__xor2_2 _21949_ (.A(_11371_),
    .B(_11568_),
    .X(_11569_));
 sky130_fd_sc_hd__buf_1 _21950_ (.A(_11569_),
    .X(_11570_));
 sky130_fd_sc_hd__buf_1 _21951_ (.A(_11570_),
    .X(_11571_));
 sky130_fd_sc_hd__xor2_2 _21952_ (.A(iY[1]),
    .B(iY[33]),
    .X(_11572_));
 sky130_fd_sc_hd__xor2_2 _21953_ (.A(_11375_),
    .B(_11572_),
    .X(_11574_));
 sky130_fd_sc_hd__buf_1 _21954_ (.A(_11574_),
    .X(_11575_));
 sky130_fd_sc_hd__buf_1 _21955_ (.A(_11575_),
    .X(_11576_));
 sky130_fd_sc_hd__nand2_2 _21956_ (.A(_11371_),
    .B(_11372_),
    .Y(_11577_));
 sky130_fd_sc_hd__buf_1 _21957_ (.A(_11577_),
    .X(_11578_));
 sky130_fd_sc_hd__buf_1 _21958_ (.A(_11578_),
    .X(_11579_));
 sky130_fd_sc_hd__o22a_2 _21959_ (.A1(_11567_),
    .A2(_11571_),
    .B1(_11576_),
    .B2(_11579_),
    .X(_11580_));
 sky130_fd_sc_hd__xnor2_2 _21960_ (.A(_11371_),
    .B(_11568_),
    .Y(_11581_));
 sky130_fd_sc_hd__xnor2_2 _21961_ (.A(_11375_),
    .B(_11572_),
    .Y(_11582_));
 sky130_fd_sc_hd__buf_4 _21962_ (.A(_11582_),
    .X(_11583_));
 sky130_fd_sc_hd__buf_4 _21963_ (.A(_11583_),
    .X(_11585_));
 sky130_fd_sc_hd__nand2_2 _21964_ (.A(_11581_),
    .B(_11585_),
    .Y(_11586_));
 sky130_fd_sc_hd__nor2_2 _21965_ (.A(_11382_),
    .B(_11586_),
    .Y(_11587_));
 sky130_fd_sc_hd__a22oi_2 _21966_ (.A1(iX[33]),
    .A2(iY[32]),
    .B1(iY[33]),
    .B2(iX[32]),
    .Y(_11588_));
 sky130_fd_sc_hd__and4_2 _21967_ (.A(iX[33]),
    .B(iX[32]),
    .C(iY[32]),
    .D(iY[33]),
    .X(_11589_));
 sky130_fd_sc_hd__nor2_2 _21968_ (.A(_11588_),
    .B(_11589_),
    .Y(_11590_));
 sky130_fd_sc_hd__o21a_2 _21969_ (.A1(_11580_),
    .A2(_11587_),
    .B1(_11590_),
    .X(_11591_));
 sky130_fd_sc_hd__nor3_2 _21970_ (.A(_11580_),
    .B(_11587_),
    .C(_11590_),
    .Y(_11592_));
 sky130_fd_sc_hd__nor2_2 _21971_ (.A(_11591_),
    .B(_11592_),
    .Y(_11593_));
 sky130_fd_sc_hd__nor2_2 _21972_ (.A(_11563_),
    .B(_11593_),
    .Y(_11594_));
 sky130_fd_sc_hd__and2_2 _21973_ (.A(_11563_),
    .B(_11593_),
    .X(_11596_));
 sky130_fd_sc_hd__nor2_2 _21974_ (.A(_11594_),
    .B(_11596_),
    .Y(_11597_));
 sky130_fd_sc_hd__xnor2_2 _21975_ (.A(oO[1]),
    .B(_11597_),
    .Y(_11598_));
 sky130_fd_sc_hd__and3_2 _21976_ (.A(_11560_),
    .B(_11561_),
    .C(_11598_),
    .X(_11599_));
 sky130_fd_sc_hd__a21o_2 _21977_ (.A1(_11560_),
    .A2(_11561_),
    .B1(_11598_),
    .X(_11600_));
 sky130_fd_sc_hd__and2b_2 _21978_ (.A_N(_11599_),
    .B(_11600_),
    .X(_11601_));
 sky130_fd_sc_hd__xor2_2 _21979_ (.A(_11386_),
    .B(_11601_),
    .X(oO[33]));
 sky130_fd_sc_hd__inv_2 _21980_ (.A(_11557_),
    .Y(_11602_));
 sky130_fd_sc_hd__nor2_2 _21981_ (.A(_11554_),
    .B(_11555_),
    .Y(_11603_));
 sky130_fd_sc_hd__and2_2 _21982_ (.A(_11495_),
    .B(_11543_),
    .X(_11604_));
 sky130_fd_sc_hd__and2_2 _21983_ (.A(_11424_),
    .B(_11445_),
    .X(_11606_));
 sky130_fd_sc_hd__and2b_2 _21984_ (.A_N(_11403_),
    .B(_11405_),
    .X(_11607_));
 sky130_fd_sc_hd__and3_2 _21985_ (.A(iY[3]),
    .B(iX[31]),
    .C(_11395_),
    .X(_11608_));
 sky130_fd_sc_hd__a21oi_2 _21986_ (.A1(iY[3]),
    .A2(iX[31]),
    .B1(_11395_),
    .Y(_11609_));
 sky130_fd_sc_hd__and4bb_2 _21987_ (.A_N(_11608_),
    .B_N(_11609_),
    .C(iY[5]),
    .D(iX[29]),
    .X(_11610_));
 sky130_fd_sc_hd__o2bb2a_2 _21988_ (.A1_N(iY[5]),
    .A2_N(iX[29]),
    .B1(_11608_),
    .B2(_11609_),
    .X(_11611_));
 sky130_fd_sc_hd__nor2_2 _21989_ (.A(_11610_),
    .B(_11611_),
    .Y(_11612_));
 sky130_fd_sc_hd__a21oi_2 _21990_ (.A1(_11394_),
    .A2(_11402_),
    .B1(_11325_),
    .Y(_11613_));
 sky130_fd_sc_hd__xnor2_2 _21991_ (.A(_11612_),
    .B(_11613_),
    .Y(_11614_));
 sky130_fd_sc_hd__o21ba_2 _21992_ (.A1(_11410_),
    .A2(_11412_),
    .B1_N(_11408_),
    .X(_11615_));
 sky130_fd_sc_hd__and3_2 _21993_ (.A(iY[3]),
    .B(iX[29]),
    .C(_11395_),
    .X(_11617_));
 sky130_fd_sc_hd__and4_2 _21994_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[27]),
    .D(iX[28]),
    .X(_11618_));
 sky130_fd_sc_hd__a22oi_2 _21995_ (.A1(iY[7]),
    .A2(iX[27]),
    .B1(iX[28]),
    .B2(iY[6]),
    .Y(_11619_));
 sky130_fd_sc_hd__and4bb_2 _21996_ (.A_N(_11618_),
    .B_N(_11619_),
    .C(iY[8]),
    .D(iX[26]),
    .X(_11620_));
 sky130_fd_sc_hd__o2bb2a_2 _21997_ (.A1_N(iY[8]),
    .A2_N(iX[26]),
    .B1(_11618_),
    .B2(_11619_),
    .X(_11621_));
 sky130_fd_sc_hd__nor2_2 _21998_ (.A(_11620_),
    .B(_11621_),
    .Y(_11622_));
 sky130_fd_sc_hd__o21ai_2 _21999_ (.A1(_11617_),
    .A2(_11401_),
    .B1(_11622_),
    .Y(_11623_));
 sky130_fd_sc_hd__or3_2 _22000_ (.A(_11617_),
    .B(_11401_),
    .C(_11622_),
    .X(_11624_));
 sky130_fd_sc_hd__and2_2 _22001_ (.A(_11623_),
    .B(_11624_),
    .X(_11625_));
 sky130_fd_sc_hd__xnor2_2 _22002_ (.A(_11615_),
    .B(_11625_),
    .Y(_11626_));
 sky130_fd_sc_hd__and2_2 _22003_ (.A(_11614_),
    .B(_11626_),
    .X(_11628_));
 sky130_fd_sc_hd__nor2_2 _22004_ (.A(_11614_),
    .B(_11626_),
    .Y(_11629_));
 sky130_fd_sc_hd__or2_2 _22005_ (.A(_11628_),
    .B(_11629_),
    .X(_11630_));
 sky130_fd_sc_hd__o21ba_2 _22006_ (.A1(_11607_),
    .A2(_11418_),
    .B1_N(_11630_),
    .X(_11631_));
 sky130_fd_sc_hd__or3b_2 _22007_ (.A(_11607_),
    .B(_11418_),
    .C_N(_11630_),
    .X(_11632_));
 sky130_fd_sc_hd__or2b_2 _22008_ (.A(_11631_),
    .B_N(_11632_),
    .X(_11633_));
 sky130_fd_sc_hd__and2b_2 _22009_ (.A_N(_11437_),
    .B(_11436_),
    .X(_11634_));
 sky130_fd_sc_hd__a21oi_2 _22010_ (.A1(_11430_),
    .A2(_11438_),
    .B1(_11634_),
    .Y(_11635_));
 sky130_fd_sc_hd__or2b_2 _22011_ (.A(_11407_),
    .B_N(_11413_),
    .X(_11636_));
 sky130_fd_sc_hd__and4_2 _22012_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[21]),
    .D(iX[22]),
    .X(_11637_));
 sky130_fd_sc_hd__a22oi_2 _22013_ (.A1(iY[13]),
    .A2(iX[21]),
    .B1(iX[22]),
    .B2(iY[12]),
    .Y(_11639_));
 sky130_fd_sc_hd__nor2_2 _22014_ (.A(_11637_),
    .B(_11639_),
    .Y(_11640_));
 sky130_fd_sc_hd__nand2_2 _22015_ (.A(iY[14]),
    .B(iX[20]),
    .Y(_11641_));
 sky130_fd_sc_hd__xnor2_2 _22016_ (.A(_11640_),
    .B(_11641_),
    .Y(_11642_));
 sky130_fd_sc_hd__and4_2 _22017_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[24]),
    .D(iX[25]),
    .X(_11643_));
 sky130_fd_sc_hd__a22oi_2 _22018_ (.A1(iY[10]),
    .A2(iX[24]),
    .B1(iX[25]),
    .B2(iY[9]),
    .Y(_11644_));
 sky130_fd_sc_hd__nor2_2 _22019_ (.A(_11643_),
    .B(_11644_),
    .Y(_11645_));
 sky130_fd_sc_hd__nand2_2 _22020_ (.A(iY[11]),
    .B(iX[23]),
    .Y(_11646_));
 sky130_fd_sc_hd__xnor2_2 _22021_ (.A(_11645_),
    .B(_11646_),
    .Y(_11647_));
 sky130_fd_sc_hd__o21ba_2 _22022_ (.A1(_11433_),
    .A2(_11435_),
    .B1_N(_11432_),
    .X(_11648_));
 sky130_fd_sc_hd__xnor2_2 _22023_ (.A(_11647_),
    .B(_11648_),
    .Y(_11650_));
 sky130_fd_sc_hd__and2_2 _22024_ (.A(_11642_),
    .B(_11650_),
    .X(_11651_));
 sky130_fd_sc_hd__nor2_2 _22025_ (.A(_11642_),
    .B(_11650_),
    .Y(_11652_));
 sky130_fd_sc_hd__or2_2 _22026_ (.A(_11651_),
    .B(_11652_),
    .X(_11653_));
 sky130_fd_sc_hd__a21o_2 _22027_ (.A1(_11636_),
    .A2(_11415_),
    .B1(_11653_),
    .X(_11654_));
 sky130_fd_sc_hd__nand3_2 _22028_ (.A(_11636_),
    .B(_11415_),
    .C(_11653_),
    .Y(_11655_));
 sky130_fd_sc_hd__nand2_2 _22029_ (.A(_11654_),
    .B(_11655_),
    .Y(_11656_));
 sky130_fd_sc_hd__xnor2_2 _22030_ (.A(_11635_),
    .B(_11656_),
    .Y(_11657_));
 sky130_fd_sc_hd__xor2_2 _22031_ (.A(_11633_),
    .B(_11657_),
    .X(_11658_));
 sky130_fd_sc_hd__o21ai_2 _22032_ (.A1(_11422_),
    .A2(_11606_),
    .B1(_11658_),
    .Y(_11659_));
 sky130_fd_sc_hd__or3_2 _22033_ (.A(_11422_),
    .B(_11606_),
    .C(_11658_),
    .X(_11661_));
 sky130_fd_sc_hd__and2_2 _22034_ (.A(_11659_),
    .B(_11661_),
    .X(_11662_));
 sky130_fd_sc_hd__and2b_2 _22035_ (.A_N(_11480_),
    .B(_11482_),
    .X(_11663_));
 sky130_fd_sc_hd__and4_2 _22036_ (.A(iX[12]),
    .B(iX[13]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_11664_));
 sky130_fd_sc_hd__a22oi_2 _22037_ (.A1(iX[13]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[12]),
    .Y(_11665_));
 sky130_fd_sc_hd__nor2_2 _22038_ (.A(_11664_),
    .B(_11665_),
    .Y(_11666_));
 sky130_fd_sc_hd__nand2_2 _22039_ (.A(iX[11]),
    .B(iY[23]),
    .Y(_11667_));
 sky130_fd_sc_hd__xnor2_2 _22040_ (.A(_11666_),
    .B(_11667_),
    .Y(_11668_));
 sky130_fd_sc_hd__and4_2 _22041_ (.A(iX[15]),
    .B(iX[16]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_11669_));
 sky130_fd_sc_hd__a22oi_2 _22042_ (.A1(iX[16]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[15]),
    .Y(_11670_));
 sky130_fd_sc_hd__nor2_2 _22043_ (.A(_11669_),
    .B(_11670_),
    .Y(_11672_));
 sky130_fd_sc_hd__nand2_2 _22044_ (.A(iX[14]),
    .B(iY[20]),
    .Y(_11673_));
 sky130_fd_sc_hd__xnor2_2 _22045_ (.A(_11672_),
    .B(_11673_),
    .Y(_11674_));
 sky130_fd_sc_hd__o21ba_2 _22046_ (.A1(_11458_),
    .A2(_11460_),
    .B1_N(_11457_),
    .X(_11675_));
 sky130_fd_sc_hd__xnor2_2 _22047_ (.A(_11674_),
    .B(_11675_),
    .Y(_11676_));
 sky130_fd_sc_hd__and2_2 _22048_ (.A(_11668_),
    .B(_11676_),
    .X(_11677_));
 sky130_fd_sc_hd__nor2_2 _22049_ (.A(_11668_),
    .B(_11676_),
    .Y(_11678_));
 sky130_fd_sc_hd__or2_2 _22050_ (.A(_11677_),
    .B(_11678_),
    .X(_11679_));
 sky130_fd_sc_hd__or3_2 _22051_ (.A(_11469_),
    .B(_11472_),
    .C(_11473_),
    .X(_11680_));
 sky130_fd_sc_hd__o21ba_2 _22052_ (.A1(_11427_),
    .A2(_11429_),
    .B1_N(_11426_),
    .X(_11681_));
 sky130_fd_sc_hd__and4_2 _22053_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[18]),
    .D(iX[19]),
    .X(_11683_));
 sky130_fd_sc_hd__a22oi_2 _22054_ (.A1(iY[16]),
    .A2(iX[18]),
    .B1(iX[19]),
    .B2(iY[15]),
    .Y(_11684_));
 sky130_fd_sc_hd__and4bb_2 _22055_ (.A_N(_11683_),
    .B_N(_11684_),
    .C(iX[17]),
    .D(iY[17]),
    .X(_11685_));
 sky130_fd_sc_hd__o2bb2a_2 _22056_ (.A1_N(iX[17]),
    .A2_N(iY[17]),
    .B1(_11683_),
    .B2(_11684_),
    .X(_11686_));
 sky130_fd_sc_hd__nor2_2 _22057_ (.A(_11685_),
    .B(_11686_),
    .Y(_11687_));
 sky130_fd_sc_hd__xnor2_2 _22058_ (.A(_11681_),
    .B(_11687_),
    .Y(_11688_));
 sky130_fd_sc_hd__o21ai_2 _22059_ (.A1(_11470_),
    .A2(_11472_),
    .B1(_11688_),
    .Y(_11689_));
 sky130_fd_sc_hd__or3_2 _22060_ (.A(_11470_),
    .B(_11472_),
    .C(_11688_),
    .X(_11690_));
 sky130_fd_sc_hd__nand2_2 _22061_ (.A(_11689_),
    .B(_11690_),
    .Y(_11691_));
 sky130_fd_sc_hd__a21oi_2 _22062_ (.A1(_11680_),
    .A2(_11477_),
    .B1(_11691_),
    .Y(_11692_));
 sky130_fd_sc_hd__and3_2 _22063_ (.A(_11680_),
    .B(_11477_),
    .C(_11691_),
    .X(_11694_));
 sky130_fd_sc_hd__or3_2 _22064_ (.A(_11679_),
    .B(_11692_),
    .C(_11694_),
    .X(_11695_));
 sky130_fd_sc_hd__o21ai_2 _22065_ (.A1(_11692_),
    .A2(_11694_),
    .B1(_11679_),
    .Y(_11696_));
 sky130_fd_sc_hd__nand2_2 _22066_ (.A(_11695_),
    .B(_11696_),
    .Y(_11697_));
 sky130_fd_sc_hd__a21oi_2 _22067_ (.A1(_11440_),
    .A2(_11443_),
    .B1(_11697_),
    .Y(_11698_));
 sky130_fd_sc_hd__and3_2 _22068_ (.A(_11440_),
    .B(_11443_),
    .C(_11697_),
    .X(_11699_));
 sky130_fd_sc_hd__nor2_2 _22069_ (.A(_11698_),
    .B(_11699_),
    .Y(_11700_));
 sky130_fd_sc_hd__xnor2_2 _22070_ (.A(_11663_),
    .B(_11700_),
    .Y(_11701_));
 sky130_fd_sc_hd__xnor2_2 _22071_ (.A(_11662_),
    .B(_11701_),
    .Y(_11702_));
 sky130_fd_sc_hd__o21ba_2 _22072_ (.A1(_11447_),
    .A2(_11490_),
    .B1_N(_11702_),
    .X(_11703_));
 sky130_fd_sc_hd__or3b_2 _22073_ (.A(_11447_),
    .B(_11490_),
    .C_N(_11702_),
    .X(_11705_));
 sky130_fd_sc_hd__or2b_2 _22074_ (.A(_11703_),
    .B_N(_11705_),
    .X(_11706_));
 sky130_fd_sc_hd__or2_2 _22075_ (.A(_11535_),
    .B(_11538_),
    .X(_11707_));
 sky130_fd_sc_hd__and2_2 _22076_ (.A(_11450_),
    .B(_11488_),
    .X(_11708_));
 sky130_fd_sc_hd__or2b_2 _22077_ (.A(_11505_),
    .B_N(_11504_),
    .X(_11709_));
 sky130_fd_sc_hd__and4_2 _22078_ (.A(iX[6]),
    .B(iX[7]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_11710_));
 sky130_fd_sc_hd__a22oi_2 _22079_ (.A1(iX[7]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[6]),
    .Y(_11711_));
 sky130_fd_sc_hd__nor2_2 _22080_ (.A(_11710_),
    .B(_11711_),
    .Y(_11712_));
 sky130_fd_sc_hd__nand2_2 _22081_ (.A(iX[5]),
    .B(iY[29]),
    .Y(_11713_));
 sky130_fd_sc_hd__xnor2_2 _22082_ (.A(_11712_),
    .B(_11713_),
    .Y(_11714_));
 sky130_fd_sc_hd__o21ba_2 _22083_ (.A1(_11501_),
    .A2(_11503_),
    .B1_N(_11500_),
    .X(_11716_));
 sky130_fd_sc_hd__xnor2_2 _22084_ (.A(_11714_),
    .B(_11716_),
    .Y(_11717_));
 sky130_fd_sc_hd__nand3_2 _22085_ (.A(iX[4]),
    .B(iY[30]),
    .C(_11717_),
    .Y(_11718_));
 sky130_fd_sc_hd__a21o_2 _22086_ (.A1(iX[4]),
    .A2(iY[30]),
    .B1(_11717_),
    .X(_11719_));
 sky130_fd_sc_hd__nand2_2 _22087_ (.A(_11718_),
    .B(_11719_),
    .Y(_11720_));
 sky130_fd_sc_hd__a21oi_2 _22088_ (.A1(_11709_),
    .A2(_11507_),
    .B1(_11720_),
    .Y(_11721_));
 sky130_fd_sc_hd__and3_2 _22089_ (.A(_11709_),
    .B(_11507_),
    .C(_11720_),
    .X(_11722_));
 sky130_fd_sc_hd__nor2_2 _22090_ (.A(_11721_),
    .B(_11722_),
    .Y(_11723_));
 sky130_fd_sc_hd__nand2_2 _22091_ (.A(iX[3]),
    .B(iY[31]),
    .Y(_11724_));
 sky130_fd_sc_hd__xnor2_2 _22092_ (.A(_11723_),
    .B(_11724_),
    .Y(_11725_));
 sky130_fd_sc_hd__and2b_2 _22093_ (.A_N(_11533_),
    .B(_11520_),
    .X(_11727_));
 sky130_fd_sc_hd__or2b_2 _22094_ (.A(_11523_),
    .B_N(_11528_),
    .X(_11728_));
 sky130_fd_sc_hd__or2b_2 _22095_ (.A(_11522_),
    .B_N(_11529_),
    .X(_11729_));
 sky130_fd_sc_hd__nand2_2 _22096_ (.A(_11728_),
    .B(_11729_),
    .Y(_11730_));
 sky130_fd_sc_hd__and2b_2 _22097_ (.A_N(_11462_),
    .B(_11461_),
    .X(_11731_));
 sky130_fd_sc_hd__o21ba_2 _22098_ (.A1(_11525_),
    .A2(_11527_),
    .B1_N(_11524_),
    .X(_11732_));
 sky130_fd_sc_hd__o21ba_2 _22099_ (.A1(_11452_),
    .A2(_11455_),
    .B1_N(_11451_),
    .X(_11733_));
 sky130_fd_sc_hd__and4_2 _22100_ (.A(iX[9]),
    .B(iX[10]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_11734_));
 sky130_fd_sc_hd__a22oi_2 _22101_ (.A1(iX[10]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[9]),
    .Y(_11735_));
 sky130_fd_sc_hd__nor2_2 _22102_ (.A(_11734_),
    .B(_11735_),
    .Y(_11736_));
 sky130_fd_sc_hd__nand2_2 _22103_ (.A(iX[8]),
    .B(iY[26]),
    .Y(_11738_));
 sky130_fd_sc_hd__xnor2_2 _22104_ (.A(_11736_),
    .B(_11738_),
    .Y(_11739_));
 sky130_fd_sc_hd__xnor2_2 _22105_ (.A(_11733_),
    .B(_11739_),
    .Y(_11740_));
 sky130_fd_sc_hd__xnor2_2 _22106_ (.A(_11732_),
    .B(_11740_),
    .Y(_11741_));
 sky130_fd_sc_hd__o21a_2 _22107_ (.A1(_11731_),
    .A2(_11465_),
    .B1(_11741_),
    .X(_11742_));
 sky130_fd_sc_hd__nor3_2 _22108_ (.A(_11731_),
    .B(_11465_),
    .C(_11741_),
    .Y(_11743_));
 sky130_fd_sc_hd__nor2_2 _22109_ (.A(_11742_),
    .B(_11743_),
    .Y(_11744_));
 sky130_fd_sc_hd__xor2_2 _22110_ (.A(_11730_),
    .B(_11744_),
    .X(_11745_));
 sky130_fd_sc_hd__o21a_2 _22111_ (.A1(_11531_),
    .A2(_11727_),
    .B1(_11745_),
    .X(_11746_));
 sky130_fd_sc_hd__inv_2 _22112_ (.A(_11746_),
    .Y(_11747_));
 sky130_fd_sc_hd__or3_2 _22113_ (.A(_11531_),
    .B(_11727_),
    .C(_11745_),
    .X(_11749_));
 sky130_fd_sc_hd__and3_2 _22114_ (.A(_11725_),
    .B(_11747_),
    .C(_11749_),
    .X(_11750_));
 sky130_fd_sc_hd__inv_2 _22115_ (.A(_11750_),
    .Y(_11751_));
 sky130_fd_sc_hd__a21o_2 _22116_ (.A1(_11747_),
    .A2(_11749_),
    .B1(_11725_),
    .X(_11752_));
 sky130_fd_sc_hd__o211a_2 _22117_ (.A1(_11485_),
    .A2(_11708_),
    .B1(_11751_),
    .C1(_11752_),
    .X(_11753_));
 sky130_fd_sc_hd__a211oi_2 _22118_ (.A1(_11751_),
    .A2(_11752_),
    .B1(_11485_),
    .C1(_11708_),
    .Y(_11754_));
 sky130_fd_sc_hd__nor2_2 _22119_ (.A(_11753_),
    .B(_11754_),
    .Y(_11755_));
 sky130_fd_sc_hd__xnor2_2 _22120_ (.A(_11707_),
    .B(_11755_),
    .Y(_11756_));
 sky130_fd_sc_hd__nor2_2 _22121_ (.A(_11706_),
    .B(_11756_),
    .Y(_11757_));
 sky130_fd_sc_hd__and2_2 _22122_ (.A(_11706_),
    .B(_11756_),
    .X(_11758_));
 sky130_fd_sc_hd__nor2_2 _22123_ (.A(_11757_),
    .B(_11758_),
    .Y(_11760_));
 sky130_fd_sc_hd__o21ai_2 _22124_ (.A1(_11493_),
    .A2(_11604_),
    .B1(_11760_),
    .Y(_11761_));
 sky130_fd_sc_hd__or3_2 _22125_ (.A(_11493_),
    .B(_11604_),
    .C(_11760_),
    .X(_11762_));
 sky130_fd_sc_hd__and2_2 _22126_ (.A(_11761_),
    .B(_11762_),
    .X(_11763_));
 sky130_fd_sc_hd__and2b_2 _22127_ (.A_N(_11496_),
    .B(_11542_),
    .X(_11764_));
 sky130_fd_sc_hd__o21ba_2 _22128_ (.A1(_11498_),
    .A2(_11541_),
    .B1_N(_11764_),
    .X(_11765_));
 sky130_fd_sc_hd__xnor2_2 _22129_ (.A(_11763_),
    .B(_11765_),
    .Y(_11766_));
 sky130_fd_sc_hd__o21ai_2 _22130_ (.A1(_11545_),
    .A2(_11548_),
    .B1(_11766_),
    .Y(_11767_));
 sky130_fd_sc_hd__or3_2 _22131_ (.A(_11545_),
    .B(_11548_),
    .C(_11766_),
    .X(_11768_));
 sky130_fd_sc_hd__and2_2 _22132_ (.A(_11767_),
    .B(_11768_),
    .X(_11769_));
 sky130_fd_sc_hd__o21ba_2 _22133_ (.A1(_11512_),
    .A2(_11514_),
    .B1_N(_11511_),
    .X(_11771_));
 sky130_fd_sc_hd__xnor2_2 _22134_ (.A(_11769_),
    .B(_11771_),
    .Y(_11772_));
 sky130_fd_sc_hd__o21ai_2 _22135_ (.A1(_11552_),
    .A2(_11603_),
    .B1(_11772_),
    .Y(_11773_));
 sky130_fd_sc_hd__or3_2 _22136_ (.A(_11552_),
    .B(_11603_),
    .C(_11772_),
    .X(_11774_));
 sky130_fd_sc_hd__and2_2 _22137_ (.A(_11773_),
    .B(_11774_),
    .X(_11775_));
 sky130_fd_sc_hd__inv_2 _22138_ (.A(_11775_),
    .Y(_11776_));
 sky130_fd_sc_hd__a21o_2 _22139_ (.A1(_11602_),
    .A2(_11560_),
    .B1(_11776_),
    .X(_11777_));
 sky130_fd_sc_hd__nand3_2 _22140_ (.A(_11602_),
    .B(_11560_),
    .C(_11776_),
    .Y(_11778_));
 sky130_fd_sc_hd__and2_2 _22141_ (.A(iX[1]),
    .B(iX[33]),
    .X(_11779_));
 sky130_fd_sc_hd__a31o_4 _22142_ (.A1(iX[0]),
    .A2(iX[32]),
    .A3(_11568_),
    .B1(_11779_),
    .X(_11780_));
 sky130_fd_sc_hd__xor2_2 _22143_ (.A(iX[2]),
    .B(iX[34]),
    .X(_11782_));
 sky130_fd_sc_hd__xor2_2 _22144_ (.A(_11780_),
    .B(_11782_),
    .X(_11783_));
 sky130_fd_sc_hd__nand2_2 _22145_ (.A(_11379_),
    .B(_11783_),
    .Y(_11784_));
 sky130_fd_sc_hd__xor2_2 _22146_ (.A(_11586_),
    .B(_11784_),
    .X(_11785_));
 sky130_fd_sc_hd__nand2_2 _22147_ (.A(iY[2]),
    .B(iY[34]),
    .Y(_11786_));
 sky130_fd_sc_hd__or2_2 _22148_ (.A(iY[2]),
    .B(iY[34]),
    .X(_11787_));
 sky130_fd_sc_hd__nand2_2 _22149_ (.A(_11786_),
    .B(_11787_),
    .Y(_11788_));
 sky130_fd_sc_hd__and2_2 _22150_ (.A(iY[1]),
    .B(iY[33]),
    .X(_11789_));
 sky130_fd_sc_hd__a31oi_4 _22151_ (.A1(iY[0]),
    .A2(iY[32]),
    .A3(_11572_),
    .B1(_11789_),
    .Y(_11790_));
 sky130_fd_sc_hd__xnor2_2 _22152_ (.A(_11788_),
    .B(_11790_),
    .Y(_11791_));
 sky130_fd_sc_hd__buf_4 _22153_ (.A(_11791_),
    .X(_11793_));
 sky130_fd_sc_hd__buf_1 _22154_ (.A(_11793_),
    .X(_11794_));
 sky130_fd_sc_hd__nor2_2 _22155_ (.A(_11578_),
    .B(_11794_),
    .Y(_11795_));
 sky130_fd_sc_hd__xnor2_2 _22156_ (.A(_11785_),
    .B(_11795_),
    .Y(_11796_));
 sky130_fd_sc_hd__nor3_2 _22157_ (.A(_11382_),
    .B(_11586_),
    .C(_11796_),
    .Y(_11797_));
 sky130_fd_sc_hd__and2b_2 _22158_ (.A_N(_11587_),
    .B(_11796_),
    .X(_11798_));
 sky130_fd_sc_hd__or2_2 _22159_ (.A(_11797_),
    .B(_11798_),
    .X(_11799_));
 sky130_fd_sc_hd__a22oi_2 _22160_ (.A1(iX[33]),
    .A2(iY[33]),
    .B1(iY[34]),
    .B2(iX[32]),
    .Y(_11800_));
 sky130_fd_sc_hd__and4_4 _22161_ (.A(iX[33]),
    .B(iX[32]),
    .C(iY[33]),
    .D(iY[34]),
    .X(_11801_));
 sky130_fd_sc_hd__and4bb_2 _22162_ (.A_N(_11800_),
    .B_N(_11801_),
    .C(iY[32]),
    .D(iX[34]),
    .X(_11802_));
 sky130_fd_sc_hd__o2bb2a_2 _22163_ (.A1_N(iY[32]),
    .A2_N(iX[34]),
    .B1(_11800_),
    .B2(_11801_),
    .X(_11804_));
 sky130_fd_sc_hd__nor2_2 _22164_ (.A(_11802_),
    .B(_11804_),
    .Y(_11805_));
 sky130_fd_sc_hd__and2_2 _22165_ (.A(_11589_),
    .B(_11805_),
    .X(_11806_));
 sky130_fd_sc_hd__nor2_2 _22166_ (.A(_11589_),
    .B(_11805_),
    .Y(_11807_));
 sky130_fd_sc_hd__nor2_2 _22167_ (.A(_11806_),
    .B(_11807_),
    .Y(_11808_));
 sky130_fd_sc_hd__or2_2 _22168_ (.A(_11799_),
    .B(_11808_),
    .X(_11809_));
 sky130_fd_sc_hd__nand2_2 _22169_ (.A(_11799_),
    .B(_11808_),
    .Y(_11810_));
 sky130_fd_sc_hd__nand2_2 _22170_ (.A(_11809_),
    .B(_11810_),
    .Y(_11811_));
 sky130_fd_sc_hd__xnor2_2 _22171_ (.A(oO[2]),
    .B(_11811_),
    .Y(_11812_));
 sky130_fd_sc_hd__nor2_2 _22172_ (.A(_11591_),
    .B(_11812_),
    .Y(_11813_));
 sky130_fd_sc_hd__and2_2 _22173_ (.A(_11591_),
    .B(_11812_),
    .X(_11815_));
 sky130_fd_sc_hd__nor2_2 _22174_ (.A(_11813_),
    .B(_11815_),
    .Y(_11816_));
 sky130_fd_sc_hd__a21oi_2 _22175_ (.A1(_10843_),
    .A2(_11597_),
    .B1(_11594_),
    .Y(_11817_));
 sky130_fd_sc_hd__xnor2_2 _22176_ (.A(_11816_),
    .B(_11817_),
    .Y(_11818_));
 sky130_fd_sc_hd__and3_2 _22177_ (.A(_11777_),
    .B(_11778_),
    .C(_11818_),
    .X(_11819_));
 sky130_fd_sc_hd__a21o_2 _22178_ (.A1(_11777_),
    .A2(_11778_),
    .B1(_11818_),
    .X(_11820_));
 sky130_fd_sc_hd__or2b_2 _22179_ (.A(_11819_),
    .B_N(_11820_),
    .X(_11821_));
 sky130_fd_sc_hd__a21o_2 _22180_ (.A1(_11386_),
    .A2(_11600_),
    .B1(_11599_),
    .X(_11822_));
 sky130_fd_sc_hd__xnor2_2 _22181_ (.A(_11821_),
    .B(_11822_),
    .Y(oO[34]));
 sky130_fd_sc_hd__xor2_2 _22182_ (.A(iX[3]),
    .B(iX[35]),
    .X(_11823_));
 sky130_fd_sc_hd__and2_2 _22183_ (.A(iX[2]),
    .B(iX[34]),
    .X(_11825_));
 sky130_fd_sc_hd__a21oi_2 _22184_ (.A1(_11780_),
    .A2(_11782_),
    .B1(_11825_),
    .Y(_11826_));
 sky130_fd_sc_hd__xor2_2 _22185_ (.A(_11823_),
    .B(_11826_),
    .X(_11827_));
 sky130_fd_sc_hd__nor3_2 _22186_ (.A(_11575_),
    .B(_11784_),
    .C(_11827_),
    .Y(_11828_));
 sky130_fd_sc_hd__xnor2_2 _22187_ (.A(_11823_),
    .B(_11826_),
    .Y(_11829_));
 sky130_fd_sc_hd__a22o_2 _22188_ (.A1(_11583_),
    .A2(_11783_),
    .B1(_11829_),
    .B2(_11379_),
    .X(_11830_));
 sky130_fd_sc_hd__and2b_2 _22189_ (.A_N(_11828_),
    .B(_11830_),
    .X(_11831_));
 sky130_fd_sc_hd__nor2_2 _22190_ (.A(_11569_),
    .B(_11791_),
    .Y(_11832_));
 sky130_fd_sc_hd__xnor2_2 _22191_ (.A(_11831_),
    .B(_11832_),
    .Y(_11833_));
 sky130_fd_sc_hd__or2_2 _22192_ (.A(_11586_),
    .B(_11784_),
    .X(_11834_));
 sky130_fd_sc_hd__a21bo_2 _22193_ (.A1(_11785_),
    .A2(_11795_),
    .B1_N(_11834_),
    .X(_11836_));
 sky130_fd_sc_hd__xor2_2 _22194_ (.A(_11833_),
    .B(_11836_),
    .X(_11837_));
 sky130_fd_sc_hd__nand2_2 _22195_ (.A(iY[3]),
    .B(iY[35]),
    .Y(_11838_));
 sky130_fd_sc_hd__or2_2 _22196_ (.A(iY[3]),
    .B(iY[35]),
    .X(_11839_));
 sky130_fd_sc_hd__nand2_2 _22197_ (.A(_11838_),
    .B(_11839_),
    .Y(_11840_));
 sky130_fd_sc_hd__o21ai_4 _22198_ (.A1(_11788_),
    .A2(_11790_),
    .B1(_11786_),
    .Y(_11841_));
 sky130_fd_sc_hd__xnor2_2 _22199_ (.A(_11840_),
    .B(_11841_),
    .Y(_11842_));
 sky130_fd_sc_hd__nand2_2 _22200_ (.A(_11373_),
    .B(_11842_),
    .Y(_11843_));
 sky130_fd_sc_hd__xor2_2 _22201_ (.A(_11837_),
    .B(_11843_),
    .X(_11844_));
 sky130_fd_sc_hd__xnor2_2 _22202_ (.A(_11797_),
    .B(_11844_),
    .Y(_11845_));
 sky130_fd_sc_hd__and4_2 _22203_ (.A(iX[33]),
    .B(iX[32]),
    .C(iY[34]),
    .D(iY[35]),
    .X(_11847_));
 sky130_fd_sc_hd__a22o_2 _22204_ (.A1(iX[33]),
    .A2(iY[34]),
    .B1(iY[35]),
    .B2(iX[32]),
    .X(_11848_));
 sky130_fd_sc_hd__and2b_2 _22205_ (.A_N(_11847_),
    .B(_11848_),
    .X(_11849_));
 sky130_fd_sc_hd__nand2_2 _22206_ (.A(iY[33]),
    .B(iX[34]),
    .Y(_11850_));
 sky130_fd_sc_hd__xnor2_2 _22207_ (.A(_11849_),
    .B(_11850_),
    .Y(_11851_));
 sky130_fd_sc_hd__xnor2_2 _22208_ (.A(_11801_),
    .B(_11851_),
    .Y(_11852_));
 sky130_fd_sc_hd__nand2_2 _22209_ (.A(iY[32]),
    .B(iX[35]),
    .Y(_11853_));
 sky130_fd_sc_hd__or2_2 _22210_ (.A(_11852_),
    .B(_11853_),
    .X(_11854_));
 sky130_fd_sc_hd__nand2_2 _22211_ (.A(_11852_),
    .B(_11853_),
    .Y(_11855_));
 sky130_fd_sc_hd__and3_2 _22212_ (.A(_11802_),
    .B(_11854_),
    .C(_11855_),
    .X(_11856_));
 sky130_fd_sc_hd__and2_2 _22213_ (.A(_11854_),
    .B(_11855_),
    .X(_11858_));
 sky130_fd_sc_hd__nor2_2 _22214_ (.A(_11802_),
    .B(_11858_),
    .Y(_11859_));
 sky130_fd_sc_hd__nor2_2 _22215_ (.A(_11856_),
    .B(_11859_),
    .Y(_11860_));
 sky130_fd_sc_hd__and2_2 _22216_ (.A(_11806_),
    .B(_11860_),
    .X(_11861_));
 sky130_fd_sc_hd__nor2_2 _22217_ (.A(_11806_),
    .B(_11860_),
    .Y(_11862_));
 sky130_fd_sc_hd__nor2_2 _22218_ (.A(_11861_),
    .B(_11862_),
    .Y(_11863_));
 sky130_fd_sc_hd__xnor2_2 _22219_ (.A(_11845_),
    .B(_11863_),
    .Y(_11864_));
 sky130_fd_sc_hd__xnor2_2 _22220_ (.A(_11093_),
    .B(_11864_),
    .Y(_11865_));
 sky130_fd_sc_hd__o21ai_2 _22221_ (.A1(oO[2]),
    .A2(_11811_),
    .B1(_11809_),
    .Y(_11866_));
 sky130_fd_sc_hd__xnor2_2 _22222_ (.A(_11865_),
    .B(_11866_),
    .Y(_11867_));
 sky130_fd_sc_hd__o21bai_2 _22223_ (.A1(_11815_),
    .A2(_11817_),
    .B1_N(_11813_),
    .Y(_11869_));
 sky130_fd_sc_hd__and2b_2 _22224_ (.A_N(_11867_),
    .B(_11869_),
    .X(_11870_));
 sky130_fd_sc_hd__and2b_2 _22225_ (.A_N(_11869_),
    .B(_11867_),
    .X(_11871_));
 sky130_fd_sc_hd__nor2_2 _22226_ (.A(_11870_),
    .B(_11871_),
    .Y(_11872_));
 sky130_fd_sc_hd__or2b_2 _22227_ (.A(_11771_),
    .B_N(_11769_),
    .X(_11873_));
 sky130_fd_sc_hd__or2b_2 _22228_ (.A(_11765_),
    .B_N(_11763_),
    .X(_11874_));
 sky130_fd_sc_hd__nand2_2 _22229_ (.A(_11662_),
    .B(_11701_),
    .Y(_11875_));
 sky130_fd_sc_hd__nor2_2 _22230_ (.A(_11633_),
    .B(_11657_),
    .Y(_11876_));
 sky130_fd_sc_hd__and2b_2 _22231_ (.A_N(_11613_),
    .B(_11612_),
    .X(_11877_));
 sky130_fd_sc_hd__a22oi_2 _22232_ (.A1(iY[5]),
    .A2(iX[30]),
    .B1(iX[31]),
    .B2(iY[4]),
    .Y(_11878_));
 sky130_fd_sc_hd__and3_2 _22233_ (.A(iY[5]),
    .B(iX[31]),
    .C(_11395_),
    .X(_11880_));
 sky130_fd_sc_hd__or2_2 _22234_ (.A(_11878_),
    .B(_11880_),
    .X(_11881_));
 sky130_fd_sc_hd__or2_2 _22235_ (.A(_11618_),
    .B(_11620_),
    .X(_11882_));
 sky130_fd_sc_hd__nand2_2 _22236_ (.A(iY[7]),
    .B(iX[28]),
    .Y(_11883_));
 sky130_fd_sc_hd__nand2_2 _22237_ (.A(iY[6]),
    .B(iX[29]),
    .Y(_11884_));
 sky130_fd_sc_hd__and4_2 _22238_ (.A(iY[6]),
    .B(iY[7]),
    .C(iX[28]),
    .D(iX[29]),
    .X(_11885_));
 sky130_fd_sc_hd__a21oi_2 _22239_ (.A1(_11883_),
    .A2(_11884_),
    .B1(_11885_),
    .Y(_11886_));
 sky130_fd_sc_hd__nand2_2 _22240_ (.A(iY[8]),
    .B(iX[27]),
    .Y(_11887_));
 sky130_fd_sc_hd__xnor2_2 _22241_ (.A(_11886_),
    .B(_11887_),
    .Y(_11888_));
 sky130_fd_sc_hd__o21ai_2 _22242_ (.A1(_11608_),
    .A2(_11610_),
    .B1(_11888_),
    .Y(_11889_));
 sky130_fd_sc_hd__or3_2 _22243_ (.A(_11608_),
    .B(_11610_),
    .C(_11888_),
    .X(_11891_));
 sky130_fd_sc_hd__and2_2 _22244_ (.A(_11889_),
    .B(_11891_),
    .X(_11892_));
 sky130_fd_sc_hd__xnor2_2 _22245_ (.A(_11882_),
    .B(_11892_),
    .Y(_11893_));
 sky130_fd_sc_hd__or2_2 _22246_ (.A(_11881_),
    .B(_11893_),
    .X(_11894_));
 sky130_fd_sc_hd__nand2_2 _22247_ (.A(_11881_),
    .B(_11893_),
    .Y(_11895_));
 sky130_fd_sc_hd__and2_2 _22248_ (.A(_11894_),
    .B(_11895_),
    .X(_11896_));
 sky130_fd_sc_hd__o21a_2 _22249_ (.A1(_11877_),
    .A2(_11628_),
    .B1(_11896_),
    .X(_11897_));
 sky130_fd_sc_hd__nor3_2 _22250_ (.A(_11877_),
    .B(_11628_),
    .C(_11896_),
    .Y(_11898_));
 sky130_fd_sc_hd__and2b_2 _22251_ (.A_N(_11648_),
    .B(_11647_),
    .X(_11899_));
 sky130_fd_sc_hd__or2b_2 _22252_ (.A(_11615_),
    .B_N(_11625_),
    .X(_11900_));
 sky130_fd_sc_hd__and4_2 _22253_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[22]),
    .D(iX[23]),
    .X(_11902_));
 sky130_fd_sc_hd__a22oi_2 _22254_ (.A1(iY[13]),
    .A2(iX[22]),
    .B1(iX[23]),
    .B2(iY[12]),
    .Y(_11903_));
 sky130_fd_sc_hd__nor2_2 _22255_ (.A(_11902_),
    .B(_11903_),
    .Y(_11904_));
 sky130_fd_sc_hd__nand2_2 _22256_ (.A(iY[14]),
    .B(iX[21]),
    .Y(_11905_));
 sky130_fd_sc_hd__xnor2_2 _22257_ (.A(_11904_),
    .B(_11905_),
    .Y(_11906_));
 sky130_fd_sc_hd__and4_2 _22258_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[25]),
    .D(iX[26]),
    .X(_11907_));
 sky130_fd_sc_hd__a22oi_2 _22259_ (.A1(iY[10]),
    .A2(iX[25]),
    .B1(iX[26]),
    .B2(iY[9]),
    .Y(_11908_));
 sky130_fd_sc_hd__nor2_2 _22260_ (.A(_11907_),
    .B(_11908_),
    .Y(_11909_));
 sky130_fd_sc_hd__nand2_2 _22261_ (.A(iY[11]),
    .B(iX[24]),
    .Y(_11910_));
 sky130_fd_sc_hd__xnor2_2 _22262_ (.A(_11909_),
    .B(_11910_),
    .Y(_11911_));
 sky130_fd_sc_hd__o21ba_2 _22263_ (.A1(_11644_),
    .A2(_11646_),
    .B1_N(_11643_),
    .X(_11913_));
 sky130_fd_sc_hd__xnor2_2 _22264_ (.A(_11911_),
    .B(_11913_),
    .Y(_11914_));
 sky130_fd_sc_hd__and2_2 _22265_ (.A(_11906_),
    .B(_11914_),
    .X(_11915_));
 sky130_fd_sc_hd__nor2_2 _22266_ (.A(_11906_),
    .B(_11914_),
    .Y(_11916_));
 sky130_fd_sc_hd__or2_2 _22267_ (.A(_11915_),
    .B(_11916_),
    .X(_11917_));
 sky130_fd_sc_hd__a21o_2 _22268_ (.A1(_11623_),
    .A2(_11900_),
    .B1(_11917_),
    .X(_11918_));
 sky130_fd_sc_hd__nand3_2 _22269_ (.A(_11623_),
    .B(_11900_),
    .C(_11917_),
    .Y(_11919_));
 sky130_fd_sc_hd__o211ai_2 _22270_ (.A1(_11899_),
    .A2(_11651_),
    .B1(_11918_),
    .C1(_11919_),
    .Y(_11920_));
 sky130_fd_sc_hd__a211o_2 _22271_ (.A1(_11918_),
    .A2(_11919_),
    .B1(_11899_),
    .C1(_11651_),
    .X(_11921_));
 sky130_fd_sc_hd__and4bb_2 _22272_ (.A_N(_11897_),
    .B_N(_11898_),
    .C(_11920_),
    .D(_11921_),
    .X(_11922_));
 sky130_fd_sc_hd__a2bb2o_2 _22273_ (.A1_N(_11897_),
    .A2_N(_11898_),
    .B1(_11920_),
    .B2(_11921_),
    .X(_11924_));
 sky130_fd_sc_hd__and2b_2 _22274_ (.A_N(_11922_),
    .B(_11924_),
    .X(_11925_));
 sky130_fd_sc_hd__o21a_2 _22275_ (.A1(_11631_),
    .A2(_11876_),
    .B1(_11925_),
    .X(_11926_));
 sky130_fd_sc_hd__nor3_2 _22276_ (.A(_11631_),
    .B(_11876_),
    .C(_11925_),
    .Y(_11927_));
 sky130_fd_sc_hd__nor2_2 _22277_ (.A(_11926_),
    .B(_11927_),
    .Y(_11928_));
 sky130_fd_sc_hd__inv_2 _22278_ (.A(_11692_),
    .Y(_11929_));
 sky130_fd_sc_hd__or2_2 _22279_ (.A(_11635_),
    .B(_11656_),
    .X(_11930_));
 sky130_fd_sc_hd__and4_2 _22280_ (.A(iX[13]),
    .B(iX[14]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_11931_));
 sky130_fd_sc_hd__a22oi_2 _22281_ (.A1(iX[14]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[13]),
    .Y(_11932_));
 sky130_fd_sc_hd__nor2_2 _22282_ (.A(_11931_),
    .B(_11932_),
    .Y(_11933_));
 sky130_fd_sc_hd__nand2_2 _22283_ (.A(iX[12]),
    .B(iY[23]),
    .Y(_11934_));
 sky130_fd_sc_hd__xnor2_2 _22284_ (.A(_11933_),
    .B(_11934_),
    .Y(_11935_));
 sky130_fd_sc_hd__and4_2 _22285_ (.A(iX[16]),
    .B(iX[17]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_11936_));
 sky130_fd_sc_hd__a22oi_2 _22286_ (.A1(iX[17]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[16]),
    .Y(_11937_));
 sky130_fd_sc_hd__nor2_2 _22287_ (.A(_11936_),
    .B(_11937_),
    .Y(_11938_));
 sky130_fd_sc_hd__nand2_2 _22288_ (.A(iX[15]),
    .B(iY[20]),
    .Y(_11939_));
 sky130_fd_sc_hd__xnor2_2 _22289_ (.A(_11938_),
    .B(_11939_),
    .Y(_11940_));
 sky130_fd_sc_hd__o21ba_2 _22290_ (.A1(_11670_),
    .A2(_11673_),
    .B1_N(_11669_),
    .X(_11941_));
 sky130_fd_sc_hd__xnor2_2 _22291_ (.A(_11940_),
    .B(_11941_),
    .Y(_11942_));
 sky130_fd_sc_hd__and2_2 _22292_ (.A(_11935_),
    .B(_11942_),
    .X(_11943_));
 sky130_fd_sc_hd__nor2_2 _22293_ (.A(_11935_),
    .B(_11942_),
    .Y(_11945_));
 sky130_fd_sc_hd__or2_2 _22294_ (.A(_11943_),
    .B(_11945_),
    .X(_11946_));
 sky130_fd_sc_hd__or3_2 _22295_ (.A(_11681_),
    .B(_11685_),
    .C(_11686_),
    .X(_11947_));
 sky130_fd_sc_hd__o21ba_2 _22296_ (.A1(_11639_),
    .A2(_11641_),
    .B1_N(_11637_),
    .X(_11948_));
 sky130_fd_sc_hd__and4_2 _22297_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[19]),
    .D(iX[20]),
    .X(_11949_));
 sky130_fd_sc_hd__a22oi_2 _22298_ (.A1(iY[16]),
    .A2(iX[19]),
    .B1(iX[20]),
    .B2(iY[15]),
    .Y(_11950_));
 sky130_fd_sc_hd__and4bb_2 _22299_ (.A_N(_11949_),
    .B_N(_11950_),
    .C(iY[17]),
    .D(iX[18]),
    .X(_11951_));
 sky130_fd_sc_hd__o2bb2a_2 _22300_ (.A1_N(iY[17]),
    .A2_N(iX[18]),
    .B1(_11949_),
    .B2(_11950_),
    .X(_11952_));
 sky130_fd_sc_hd__nor2_2 _22301_ (.A(_11951_),
    .B(_11952_),
    .Y(_11953_));
 sky130_fd_sc_hd__xnor2_2 _22302_ (.A(_11948_),
    .B(_11953_),
    .Y(_11954_));
 sky130_fd_sc_hd__o21ai_2 _22303_ (.A1(_11683_),
    .A2(_11685_),
    .B1(_11954_),
    .Y(_11956_));
 sky130_fd_sc_hd__or3_2 _22304_ (.A(_11683_),
    .B(_11685_),
    .C(_11954_),
    .X(_11957_));
 sky130_fd_sc_hd__nand2_2 _22305_ (.A(_11956_),
    .B(_11957_),
    .Y(_11958_));
 sky130_fd_sc_hd__a21oi_2 _22306_ (.A1(_11947_),
    .A2(_11689_),
    .B1(_11958_),
    .Y(_11959_));
 sky130_fd_sc_hd__and3_2 _22307_ (.A(_11947_),
    .B(_11689_),
    .C(_11958_),
    .X(_11960_));
 sky130_fd_sc_hd__or3_2 _22308_ (.A(_11946_),
    .B(_11959_),
    .C(_11960_),
    .X(_11961_));
 sky130_fd_sc_hd__o21ai_2 _22309_ (.A1(_11959_),
    .A2(_11960_),
    .B1(_11946_),
    .Y(_11962_));
 sky130_fd_sc_hd__nand2_2 _22310_ (.A(_11961_),
    .B(_11962_),
    .Y(_11963_));
 sky130_fd_sc_hd__a21oi_2 _22311_ (.A1(_11654_),
    .A2(_11930_),
    .B1(_11963_),
    .Y(_11964_));
 sky130_fd_sc_hd__and3_2 _22312_ (.A(_11654_),
    .B(_11930_),
    .C(_11963_),
    .X(_11965_));
 sky130_fd_sc_hd__a211oi_2 _22313_ (.A1(_11929_),
    .A2(_11695_),
    .B1(_11964_),
    .C1(_11965_),
    .Y(_11967_));
 sky130_fd_sc_hd__o211a_2 _22314_ (.A1(_11964_),
    .A2(_11965_),
    .B1(_11929_),
    .C1(_11695_),
    .X(_11968_));
 sky130_fd_sc_hd__nor2_2 _22315_ (.A(_11967_),
    .B(_11968_),
    .Y(_11969_));
 sky130_fd_sc_hd__xnor2_2 _22316_ (.A(_11928_),
    .B(_11969_),
    .Y(_11970_));
 sky130_fd_sc_hd__a21oi_2 _22317_ (.A1(_11659_),
    .A2(_11875_),
    .B1(_11970_),
    .Y(_11971_));
 sky130_fd_sc_hd__nand3_2 _22318_ (.A(_11659_),
    .B(_11875_),
    .C(_11970_),
    .Y(_11972_));
 sky130_fd_sc_hd__and2b_2 _22319_ (.A_N(_11971_),
    .B(_11972_),
    .X(_11973_));
 sky130_fd_sc_hd__or2_2 _22320_ (.A(_11746_),
    .B(_11750_),
    .X(_11974_));
 sky130_fd_sc_hd__o21ba_2 _22321_ (.A1(_11663_),
    .A2(_11699_),
    .B1_N(_11698_),
    .X(_11975_));
 sky130_fd_sc_hd__or2b_2 _22322_ (.A(_11716_),
    .B_N(_11714_),
    .X(_11976_));
 sky130_fd_sc_hd__and4_2 _22323_ (.A(iX[7]),
    .B(iX[8]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_11978_));
 sky130_fd_sc_hd__a22oi_2 _22324_ (.A1(iX[8]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[7]),
    .Y(_11979_));
 sky130_fd_sc_hd__nor2_2 _22325_ (.A(_11978_),
    .B(_11979_),
    .Y(_11980_));
 sky130_fd_sc_hd__nand2_2 _22326_ (.A(iX[6]),
    .B(iY[29]),
    .Y(_11981_));
 sky130_fd_sc_hd__xnor2_2 _22327_ (.A(_11980_),
    .B(_11981_),
    .Y(_11982_));
 sky130_fd_sc_hd__o21ba_2 _22328_ (.A1(_11711_),
    .A2(_11713_),
    .B1_N(_11710_),
    .X(_11983_));
 sky130_fd_sc_hd__xnor2_2 _22329_ (.A(_11982_),
    .B(_11983_),
    .Y(_11984_));
 sky130_fd_sc_hd__nand3_2 _22330_ (.A(iX[5]),
    .B(iY[30]),
    .C(_11984_),
    .Y(_11985_));
 sky130_fd_sc_hd__a21o_2 _22331_ (.A1(iX[5]),
    .A2(iY[30]),
    .B1(_11984_),
    .X(_11986_));
 sky130_fd_sc_hd__nand2_2 _22332_ (.A(_11985_),
    .B(_11986_),
    .Y(_11987_));
 sky130_fd_sc_hd__a21oi_2 _22333_ (.A1(_11976_),
    .A2(_11718_),
    .B1(_11987_),
    .Y(_11989_));
 sky130_fd_sc_hd__and3_2 _22334_ (.A(_11976_),
    .B(_11718_),
    .C(_11987_),
    .X(_11990_));
 sky130_fd_sc_hd__nor2_2 _22335_ (.A(_11989_),
    .B(_11990_),
    .Y(_11991_));
 sky130_fd_sc_hd__nand2_2 _22336_ (.A(iX[4]),
    .B(iY[31]),
    .Y(_11992_));
 sky130_fd_sc_hd__xnor2_2 _22337_ (.A(_11991_),
    .B(_11992_),
    .Y(_11993_));
 sky130_fd_sc_hd__or2b_2 _22338_ (.A(_11733_),
    .B_N(_11739_),
    .X(_11994_));
 sky130_fd_sc_hd__or2b_2 _22339_ (.A(_11732_),
    .B_N(_11740_),
    .X(_11995_));
 sky130_fd_sc_hd__and2b_2 _22340_ (.A_N(_11675_),
    .B(_11674_),
    .X(_11996_));
 sky130_fd_sc_hd__o21ba_2 _22341_ (.A1(_11735_),
    .A2(_11738_),
    .B1_N(_11734_),
    .X(_11997_));
 sky130_fd_sc_hd__o21ba_2 _22342_ (.A1(_11665_),
    .A2(_11667_),
    .B1_N(_11664_),
    .X(_11998_));
 sky130_fd_sc_hd__and4_2 _22343_ (.A(iX[10]),
    .B(iX[11]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_12000_));
 sky130_fd_sc_hd__a22oi_2 _22344_ (.A1(iX[11]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[10]),
    .Y(_12001_));
 sky130_fd_sc_hd__nor2_2 _22345_ (.A(_12000_),
    .B(_12001_),
    .Y(_12002_));
 sky130_fd_sc_hd__nand2_2 _22346_ (.A(iX[9]),
    .B(iY[26]),
    .Y(_12003_));
 sky130_fd_sc_hd__xnor2_2 _22347_ (.A(_12002_),
    .B(_12003_),
    .Y(_12004_));
 sky130_fd_sc_hd__xnor2_2 _22348_ (.A(_11998_),
    .B(_12004_),
    .Y(_12005_));
 sky130_fd_sc_hd__xnor2_2 _22349_ (.A(_11997_),
    .B(_12005_),
    .Y(_12006_));
 sky130_fd_sc_hd__o21a_2 _22350_ (.A1(_11996_),
    .A2(_11677_),
    .B1(_12006_),
    .X(_12007_));
 sky130_fd_sc_hd__nor3_2 _22351_ (.A(_11996_),
    .B(_11677_),
    .C(_12006_),
    .Y(_12008_));
 sky130_fd_sc_hd__a211oi_2 _22352_ (.A1(_11994_),
    .A2(_11995_),
    .B1(_12007_),
    .C1(_12008_),
    .Y(_12009_));
 sky130_fd_sc_hd__o211a_2 _22353_ (.A1(_12007_),
    .A2(_12008_),
    .B1(_11994_),
    .C1(_11995_),
    .X(_12011_));
 sky130_fd_sc_hd__a21oi_2 _22354_ (.A1(_11730_),
    .A2(_11744_),
    .B1(_11742_),
    .Y(_12012_));
 sky130_fd_sc_hd__or3_2 _22355_ (.A(_12009_),
    .B(_12011_),
    .C(_12012_),
    .X(_12013_));
 sky130_fd_sc_hd__o21ai_2 _22356_ (.A1(_12009_),
    .A2(_12011_),
    .B1(_12012_),
    .Y(_12014_));
 sky130_fd_sc_hd__and3_2 _22357_ (.A(_11993_),
    .B(_12013_),
    .C(_12014_),
    .X(_12015_));
 sky130_fd_sc_hd__a21oi_2 _22358_ (.A1(_12013_),
    .A2(_12014_),
    .B1(_11993_),
    .Y(_12016_));
 sky130_fd_sc_hd__or3_2 _22359_ (.A(_11975_),
    .B(_12015_),
    .C(_12016_),
    .X(_12017_));
 sky130_fd_sc_hd__o21ai_2 _22360_ (.A1(_12015_),
    .A2(_12016_),
    .B1(_11975_),
    .Y(_12018_));
 sky130_fd_sc_hd__nand2_2 _22361_ (.A(_12017_),
    .B(_12018_),
    .Y(_12019_));
 sky130_fd_sc_hd__xnor2_2 _22362_ (.A(_11974_),
    .B(_12019_),
    .Y(_12020_));
 sky130_fd_sc_hd__xor2_2 _22363_ (.A(_11973_),
    .B(_12020_),
    .X(_12022_));
 sky130_fd_sc_hd__o21ai_2 _22364_ (.A1(_11703_),
    .A2(_11757_),
    .B1(_12022_),
    .Y(_12023_));
 sky130_fd_sc_hd__or3_2 _22365_ (.A(_11703_),
    .B(_11757_),
    .C(_12022_),
    .X(_12024_));
 sky130_fd_sc_hd__and2_2 _22366_ (.A(_12023_),
    .B(_12024_),
    .X(_12025_));
 sky130_fd_sc_hd__a21o_2 _22367_ (.A1(_11707_),
    .A2(_11755_),
    .B1(_11753_),
    .X(_12026_));
 sky130_fd_sc_hd__xnor2_2 _22368_ (.A(_12025_),
    .B(_12026_),
    .Y(_12027_));
 sky130_fd_sc_hd__a21o_2 _22369_ (.A1(_11761_),
    .A2(_11874_),
    .B1(_12027_),
    .X(_12028_));
 sky130_fd_sc_hd__nand3_2 _22370_ (.A(_11761_),
    .B(_11874_),
    .C(_12027_),
    .Y(_12029_));
 sky130_fd_sc_hd__and2_2 _22371_ (.A(_12028_),
    .B(_12029_),
    .X(_12030_));
 sky130_fd_sc_hd__a31o_2 _22372_ (.A1(iX[3]),
    .A2(iY[31]),
    .A3(_11723_),
    .B1(_11721_),
    .X(_12031_));
 sky130_fd_sc_hd__xnor2_2 _22373_ (.A(_12030_),
    .B(_12031_),
    .Y(_12033_));
 sky130_fd_sc_hd__a21oi_2 _22374_ (.A1(_11767_),
    .A2(_11873_),
    .B1(_12033_),
    .Y(_12034_));
 sky130_fd_sc_hd__and3_2 _22375_ (.A(_11767_),
    .B(_11873_),
    .C(_12033_),
    .X(_12035_));
 sky130_fd_sc_hd__nor2_2 _22376_ (.A(_12034_),
    .B(_12035_),
    .Y(_12036_));
 sky130_fd_sc_hd__inv_2 _22377_ (.A(_12036_),
    .Y(_12037_));
 sky130_fd_sc_hd__a21o_2 _22378_ (.A1(_11773_),
    .A2(_11777_),
    .B1(_12037_),
    .X(_12038_));
 sky130_fd_sc_hd__nand3_2 _22379_ (.A(_11773_),
    .B(_11777_),
    .C(_12037_),
    .Y(_12039_));
 sky130_fd_sc_hd__and3_2 _22380_ (.A(_11872_),
    .B(_12038_),
    .C(_12039_),
    .X(_12040_));
 sky130_fd_sc_hd__a21oi_2 _22381_ (.A1(_12038_),
    .A2(_12039_),
    .B1(_11872_),
    .Y(_12041_));
 sky130_fd_sc_hd__nor2_2 _22382_ (.A(_12040_),
    .B(_12041_),
    .Y(_12042_));
 sky130_fd_sc_hd__a21oi_2 _22383_ (.A1(_11820_),
    .A2(_11822_),
    .B1(_11819_),
    .Y(_12044_));
 sky130_fd_sc_hd__xnor2_2 _22384_ (.A(_12042_),
    .B(_12044_),
    .Y(oO[35]));
 sky130_fd_sc_hd__nand2_2 _22385_ (.A(_12030_),
    .B(_12031_),
    .Y(_12045_));
 sky130_fd_sc_hd__nand2_2 _22386_ (.A(_12025_),
    .B(_12026_),
    .Y(_12046_));
 sky130_fd_sc_hd__and2_2 _22387_ (.A(_11928_),
    .B(_11969_),
    .X(_12047_));
 sky130_fd_sc_hd__nand2_2 _22388_ (.A(iY[5]),
    .B(iX[31]),
    .Y(_12048_));
 sky130_fd_sc_hd__a31o_2 _22389_ (.A1(iY[8]),
    .A2(iX[27]),
    .A3(_11886_),
    .B1(_11885_),
    .X(_12049_));
 sky130_fd_sc_hd__nand2_2 _22390_ (.A(iY[7]),
    .B(iX[30]),
    .Y(_12050_));
 sky130_fd_sc_hd__nor2_2 _22391_ (.A(_11884_),
    .B(_12050_),
    .Y(_12051_));
 sky130_fd_sc_hd__nand2_2 _22392_ (.A(iY[6]),
    .B(iX[30]),
    .Y(_12052_));
 sky130_fd_sc_hd__a21boi_2 _22393_ (.A1(iY[7]),
    .A2(iX[29]),
    .B1_N(_12052_),
    .Y(_12054_));
 sky130_fd_sc_hd__and4bb_2 _22394_ (.A_N(_12051_),
    .B_N(_12054_),
    .C(iY[8]),
    .D(iX[28]),
    .X(_12055_));
 sky130_fd_sc_hd__o2bb2a_2 _22395_ (.A1_N(iY[8]),
    .A2_N(iX[28]),
    .B1(_12051_),
    .B2(_12054_),
    .X(_12056_));
 sky130_fd_sc_hd__nor2_2 _22396_ (.A(_12055_),
    .B(_12056_),
    .Y(_12057_));
 sky130_fd_sc_hd__nand2_2 _22397_ (.A(_11880_),
    .B(_12057_),
    .Y(_12058_));
 sky130_fd_sc_hd__or2_2 _22398_ (.A(_11880_),
    .B(_12057_),
    .X(_12059_));
 sky130_fd_sc_hd__nand2_2 _22399_ (.A(_12058_),
    .B(_12059_),
    .Y(_12060_));
 sky130_fd_sc_hd__xor2_2 _22400_ (.A(_12049_),
    .B(_12060_),
    .X(_12061_));
 sky130_fd_sc_hd__or2_2 _22401_ (.A(_12048_),
    .B(_12061_),
    .X(_12062_));
 sky130_fd_sc_hd__nand2_2 _22402_ (.A(_12048_),
    .B(_12061_),
    .Y(_12063_));
 sky130_fd_sc_hd__and2_2 _22403_ (.A(_12062_),
    .B(_12063_),
    .X(_12065_));
 sky130_fd_sc_hd__xnor2_2 _22404_ (.A(_11894_),
    .B(_12065_),
    .Y(_12066_));
 sky130_fd_sc_hd__and2b_2 _22405_ (.A_N(_11913_),
    .B(_11911_),
    .X(_12067_));
 sky130_fd_sc_hd__nand2_2 _22406_ (.A(_11882_),
    .B(_11892_),
    .Y(_12068_));
 sky130_fd_sc_hd__and4_2 _22407_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[23]),
    .D(iX[24]),
    .X(_12069_));
 sky130_fd_sc_hd__a22oi_2 _22408_ (.A1(iY[13]),
    .A2(iX[23]),
    .B1(iX[24]),
    .B2(iY[12]),
    .Y(_12070_));
 sky130_fd_sc_hd__nor2_2 _22409_ (.A(_12069_),
    .B(_12070_),
    .Y(_12071_));
 sky130_fd_sc_hd__nand2_2 _22410_ (.A(iY[14]),
    .B(iX[22]),
    .Y(_12072_));
 sky130_fd_sc_hd__xnor2_2 _22411_ (.A(_12071_),
    .B(_12072_),
    .Y(_12073_));
 sky130_fd_sc_hd__and4_2 _22412_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[26]),
    .D(iX[27]),
    .X(_12074_));
 sky130_fd_sc_hd__a22oi_2 _22413_ (.A1(iY[10]),
    .A2(iX[26]),
    .B1(iX[27]),
    .B2(iY[9]),
    .Y(_12076_));
 sky130_fd_sc_hd__nor2_2 _22414_ (.A(_12074_),
    .B(_12076_),
    .Y(_12077_));
 sky130_fd_sc_hd__nand2_2 _22415_ (.A(iY[11]),
    .B(iX[25]),
    .Y(_12078_));
 sky130_fd_sc_hd__xnor2_2 _22416_ (.A(_12077_),
    .B(_12078_),
    .Y(_12079_));
 sky130_fd_sc_hd__o21ba_2 _22417_ (.A1(_11908_),
    .A2(_11910_),
    .B1_N(_11907_),
    .X(_12080_));
 sky130_fd_sc_hd__xnor2_2 _22418_ (.A(_12079_),
    .B(_12080_),
    .Y(_12081_));
 sky130_fd_sc_hd__and2_2 _22419_ (.A(_12073_),
    .B(_12081_),
    .X(_12082_));
 sky130_fd_sc_hd__nor2_2 _22420_ (.A(_12073_),
    .B(_12081_),
    .Y(_12083_));
 sky130_fd_sc_hd__or2_2 _22421_ (.A(_12082_),
    .B(_12083_),
    .X(_12084_));
 sky130_fd_sc_hd__a21o_2 _22422_ (.A1(_11889_),
    .A2(_12068_),
    .B1(_12084_),
    .X(_12085_));
 sky130_fd_sc_hd__nand3_2 _22423_ (.A(_11889_),
    .B(_12068_),
    .C(_12084_),
    .Y(_12087_));
 sky130_fd_sc_hd__o211ai_2 _22424_ (.A1(_12067_),
    .A2(_11915_),
    .B1(_12085_),
    .C1(_12087_),
    .Y(_12088_));
 sky130_fd_sc_hd__a211o_2 _22425_ (.A1(_12085_),
    .A2(_12087_),
    .B1(_12067_),
    .C1(_11915_),
    .X(_12089_));
 sky130_fd_sc_hd__nand3_2 _22426_ (.A(_12066_),
    .B(_12088_),
    .C(_12089_),
    .Y(_12090_));
 sky130_fd_sc_hd__a21o_2 _22427_ (.A1(_12088_),
    .A2(_12089_),
    .B1(_12066_),
    .X(_12091_));
 sky130_fd_sc_hd__o211a_2 _22428_ (.A1(_11897_),
    .A2(_11922_),
    .B1(_12090_),
    .C1(_12091_),
    .X(_12092_));
 sky130_fd_sc_hd__a211oi_2 _22429_ (.A1(_12090_),
    .A2(_12091_),
    .B1(_11897_),
    .C1(_11922_),
    .Y(_12093_));
 sky130_fd_sc_hd__inv_2 _22430_ (.A(_11959_),
    .Y(_12094_));
 sky130_fd_sc_hd__and4_2 _22431_ (.A(iX[14]),
    .B(iX[15]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_12095_));
 sky130_fd_sc_hd__a22oi_2 _22432_ (.A1(iX[15]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[14]),
    .Y(_12096_));
 sky130_fd_sc_hd__nor2_2 _22433_ (.A(_12095_),
    .B(_12096_),
    .Y(_12098_));
 sky130_fd_sc_hd__nand2_2 _22434_ (.A(iX[13]),
    .B(iY[23]),
    .Y(_12099_));
 sky130_fd_sc_hd__xnor2_2 _22435_ (.A(_12098_),
    .B(_12099_),
    .Y(_12100_));
 sky130_fd_sc_hd__and4_2 _22436_ (.A(iX[17]),
    .B(iX[18]),
    .C(iY[18]),
    .D(iY[19]),
    .X(_12101_));
 sky130_fd_sc_hd__a22oi_2 _22437_ (.A1(iX[18]),
    .A2(iY[18]),
    .B1(iY[19]),
    .B2(iX[17]),
    .Y(_12102_));
 sky130_fd_sc_hd__nor2_2 _22438_ (.A(_12101_),
    .B(_12102_),
    .Y(_12103_));
 sky130_fd_sc_hd__nand2_2 _22439_ (.A(iX[16]),
    .B(iY[20]),
    .Y(_12104_));
 sky130_fd_sc_hd__xnor2_2 _22440_ (.A(_12103_),
    .B(_12104_),
    .Y(_12105_));
 sky130_fd_sc_hd__o21ba_2 _22441_ (.A1(_11937_),
    .A2(_11939_),
    .B1_N(_11936_),
    .X(_12106_));
 sky130_fd_sc_hd__xnor2_2 _22442_ (.A(_12105_),
    .B(_12106_),
    .Y(_12107_));
 sky130_fd_sc_hd__and2_2 _22443_ (.A(_12100_),
    .B(_12107_),
    .X(_12109_));
 sky130_fd_sc_hd__nor2_2 _22444_ (.A(_12100_),
    .B(_12107_),
    .Y(_12110_));
 sky130_fd_sc_hd__or2_2 _22445_ (.A(_12109_),
    .B(_12110_),
    .X(_12111_));
 sky130_fd_sc_hd__or3_2 _22446_ (.A(_11948_),
    .B(_11951_),
    .C(_11952_),
    .X(_12112_));
 sky130_fd_sc_hd__o21ba_2 _22447_ (.A1(_11903_),
    .A2(_11905_),
    .B1_N(_11902_),
    .X(_12113_));
 sky130_fd_sc_hd__and4_2 _22448_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[20]),
    .D(iX[21]),
    .X(_12114_));
 sky130_fd_sc_hd__a22oi_2 _22449_ (.A1(iY[16]),
    .A2(iX[20]),
    .B1(iX[21]),
    .B2(iY[15]),
    .Y(_12115_));
 sky130_fd_sc_hd__and4bb_2 _22450_ (.A_N(_12114_),
    .B_N(_12115_),
    .C(iY[17]),
    .D(iX[19]),
    .X(_12116_));
 sky130_fd_sc_hd__o2bb2a_2 _22451_ (.A1_N(iY[17]),
    .A2_N(iX[19]),
    .B1(_12114_),
    .B2(_12115_),
    .X(_12117_));
 sky130_fd_sc_hd__nor2_2 _22452_ (.A(_12116_),
    .B(_12117_),
    .Y(_12118_));
 sky130_fd_sc_hd__xnor2_2 _22453_ (.A(_12113_),
    .B(_12118_),
    .Y(_12120_));
 sky130_fd_sc_hd__o21ai_2 _22454_ (.A1(_11949_),
    .A2(_11951_),
    .B1(_12120_),
    .Y(_12121_));
 sky130_fd_sc_hd__or3_2 _22455_ (.A(_11949_),
    .B(_11951_),
    .C(_12120_),
    .X(_12122_));
 sky130_fd_sc_hd__nand2_2 _22456_ (.A(_12121_),
    .B(_12122_),
    .Y(_12123_));
 sky130_fd_sc_hd__a21oi_2 _22457_ (.A1(_12112_),
    .A2(_11956_),
    .B1(_12123_),
    .Y(_12124_));
 sky130_fd_sc_hd__and3_2 _22458_ (.A(_12112_),
    .B(_11956_),
    .C(_12123_),
    .X(_12125_));
 sky130_fd_sc_hd__or3_2 _22459_ (.A(_12111_),
    .B(_12124_),
    .C(_12125_),
    .X(_12126_));
 sky130_fd_sc_hd__o21ai_2 _22460_ (.A1(_12124_),
    .A2(_12125_),
    .B1(_12111_),
    .Y(_12127_));
 sky130_fd_sc_hd__nand2_2 _22461_ (.A(_12126_),
    .B(_12127_),
    .Y(_12128_));
 sky130_fd_sc_hd__a21oi_2 _22462_ (.A1(_11918_),
    .A2(_11920_),
    .B1(_12128_),
    .Y(_12129_));
 sky130_fd_sc_hd__and3_2 _22463_ (.A(_11918_),
    .B(_11920_),
    .C(_12128_),
    .X(_12131_));
 sky130_fd_sc_hd__a211oi_2 _22464_ (.A1(_12094_),
    .A2(_11961_),
    .B1(_12129_),
    .C1(_12131_),
    .Y(_12132_));
 sky130_fd_sc_hd__o211a_2 _22465_ (.A1(_12129_),
    .A2(_12131_),
    .B1(_12094_),
    .C1(_11961_),
    .X(_12133_));
 sky130_fd_sc_hd__nor4_2 _22466_ (.A(_12092_),
    .B(_12093_),
    .C(_12132_),
    .D(_12133_),
    .Y(_12134_));
 sky130_fd_sc_hd__o22a_2 _22467_ (.A1(_12092_),
    .A2(_12093_),
    .B1(_12132_),
    .B2(_12133_),
    .X(_12135_));
 sky130_fd_sc_hd__nor2_2 _22468_ (.A(_12134_),
    .B(_12135_),
    .Y(_12136_));
 sky130_fd_sc_hd__o21a_2 _22469_ (.A1(_11926_),
    .A2(_12047_),
    .B1(_12136_),
    .X(_12137_));
 sky130_fd_sc_hd__nor3_2 _22470_ (.A(_11926_),
    .B(_12047_),
    .C(_12136_),
    .Y(_12138_));
 sky130_fd_sc_hd__nor2_2 _22471_ (.A(_12137_),
    .B(_12138_),
    .Y(_12139_));
 sky130_fd_sc_hd__inv_2 _22472_ (.A(_12013_),
    .Y(_12140_));
 sky130_fd_sc_hd__nor2_2 _22473_ (.A(_12140_),
    .B(_12015_),
    .Y(_12142_));
 sky130_fd_sc_hd__or2b_2 _22474_ (.A(_11983_),
    .B_N(_11982_),
    .X(_12143_));
 sky130_fd_sc_hd__and4_2 _22475_ (.A(iX[8]),
    .B(iX[9]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_12144_));
 sky130_fd_sc_hd__a22oi_2 _22476_ (.A1(iX[9]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[8]),
    .Y(_12145_));
 sky130_fd_sc_hd__nor2_2 _22477_ (.A(_12144_),
    .B(_12145_),
    .Y(_12146_));
 sky130_fd_sc_hd__nand2_2 _22478_ (.A(iX[7]),
    .B(iY[29]),
    .Y(_12147_));
 sky130_fd_sc_hd__xnor2_2 _22479_ (.A(_12146_),
    .B(_12147_),
    .Y(_12148_));
 sky130_fd_sc_hd__o21ba_2 _22480_ (.A1(_11979_),
    .A2(_11981_),
    .B1_N(_11978_),
    .X(_12149_));
 sky130_fd_sc_hd__xnor2_2 _22481_ (.A(_12148_),
    .B(_12149_),
    .Y(_12150_));
 sky130_fd_sc_hd__nand3_2 _22482_ (.A(iX[6]),
    .B(iY[30]),
    .C(_12150_),
    .Y(_12151_));
 sky130_fd_sc_hd__a21o_2 _22483_ (.A1(iX[6]),
    .A2(iY[30]),
    .B1(_12150_),
    .X(_12153_));
 sky130_fd_sc_hd__nand2_2 _22484_ (.A(_12151_),
    .B(_12153_),
    .Y(_12154_));
 sky130_fd_sc_hd__a21oi_2 _22485_ (.A1(_12143_),
    .A2(_11985_),
    .B1(_12154_),
    .Y(_12155_));
 sky130_fd_sc_hd__and3_2 _22486_ (.A(_12143_),
    .B(_11985_),
    .C(_12154_),
    .X(_12156_));
 sky130_fd_sc_hd__nor2_2 _22487_ (.A(_12155_),
    .B(_12156_),
    .Y(_12157_));
 sky130_fd_sc_hd__nand2_2 _22488_ (.A(iX[5]),
    .B(iY[31]),
    .Y(_12158_));
 sky130_fd_sc_hd__xnor2_2 _22489_ (.A(_12157_),
    .B(_12158_),
    .Y(_12159_));
 sky130_fd_sc_hd__or2b_2 _22490_ (.A(_11998_),
    .B_N(_12004_),
    .X(_12160_));
 sky130_fd_sc_hd__or2b_2 _22491_ (.A(_11997_),
    .B_N(_12005_),
    .X(_12161_));
 sky130_fd_sc_hd__and2b_2 _22492_ (.A_N(_11941_),
    .B(_11940_),
    .X(_12162_));
 sky130_fd_sc_hd__o21ba_2 _22493_ (.A1(_12001_),
    .A2(_12003_),
    .B1_N(_12000_),
    .X(_12164_));
 sky130_fd_sc_hd__o21ba_2 _22494_ (.A1(_11932_),
    .A2(_11934_),
    .B1_N(_11931_),
    .X(_12165_));
 sky130_fd_sc_hd__and4_2 _22495_ (.A(iX[11]),
    .B(iX[12]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_12166_));
 sky130_fd_sc_hd__a22oi_2 _22496_ (.A1(iX[12]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[11]),
    .Y(_12167_));
 sky130_fd_sc_hd__nor2_2 _22497_ (.A(_12166_),
    .B(_12167_),
    .Y(_12168_));
 sky130_fd_sc_hd__nand2_2 _22498_ (.A(iX[10]),
    .B(iY[26]),
    .Y(_12169_));
 sky130_fd_sc_hd__xnor2_2 _22499_ (.A(_12168_),
    .B(_12169_),
    .Y(_12170_));
 sky130_fd_sc_hd__xnor2_2 _22500_ (.A(_12165_),
    .B(_12170_),
    .Y(_12171_));
 sky130_fd_sc_hd__xnor2_2 _22501_ (.A(_12164_),
    .B(_12171_),
    .Y(_12172_));
 sky130_fd_sc_hd__o21a_2 _22502_ (.A1(_12162_),
    .A2(_11943_),
    .B1(_12172_),
    .X(_12173_));
 sky130_fd_sc_hd__nor3_2 _22503_ (.A(_12162_),
    .B(_11943_),
    .C(_12172_),
    .Y(_12175_));
 sky130_fd_sc_hd__a211oi_2 _22504_ (.A1(_12160_),
    .A2(_12161_),
    .B1(_12173_),
    .C1(_12175_),
    .Y(_12176_));
 sky130_fd_sc_hd__o211a_2 _22505_ (.A1(_12173_),
    .A2(_12175_),
    .B1(_12160_),
    .C1(_12161_),
    .X(_12177_));
 sky130_fd_sc_hd__nor2_2 _22506_ (.A(_12007_),
    .B(_12009_),
    .Y(_12178_));
 sky130_fd_sc_hd__or3_2 _22507_ (.A(_12176_),
    .B(_12177_),
    .C(_12178_),
    .X(_12179_));
 sky130_fd_sc_hd__o21ai_2 _22508_ (.A1(_12176_),
    .A2(_12177_),
    .B1(_12178_),
    .Y(_12180_));
 sky130_fd_sc_hd__and3_2 _22509_ (.A(_12159_),
    .B(_12179_),
    .C(_12180_),
    .X(_12181_));
 sky130_fd_sc_hd__a21oi_2 _22510_ (.A1(_12179_),
    .A2(_12180_),
    .B1(_12159_),
    .Y(_12182_));
 sky130_fd_sc_hd__nor2_2 _22511_ (.A(_12181_),
    .B(_12182_),
    .Y(_12183_));
 sky130_fd_sc_hd__o21a_2 _22512_ (.A1(_11964_),
    .A2(_11967_),
    .B1(_12183_),
    .X(_12184_));
 sky130_fd_sc_hd__nor3_2 _22513_ (.A(_11964_),
    .B(_11967_),
    .C(_12183_),
    .Y(_12186_));
 sky130_fd_sc_hd__nor2_2 _22514_ (.A(_12184_),
    .B(_12186_),
    .Y(_12187_));
 sky130_fd_sc_hd__xnor2_2 _22515_ (.A(_12142_),
    .B(_12187_),
    .Y(_12188_));
 sky130_fd_sc_hd__xnor2_2 _22516_ (.A(_12139_),
    .B(_12188_),
    .Y(_12189_));
 sky130_fd_sc_hd__a21oi_2 _22517_ (.A1(_11972_),
    .A2(_12020_),
    .B1(_11971_),
    .Y(_12190_));
 sky130_fd_sc_hd__xnor2_2 _22518_ (.A(_12189_),
    .B(_12190_),
    .Y(_12191_));
 sky130_fd_sc_hd__a21bo_2 _22519_ (.A1(_11974_),
    .A2(_12018_),
    .B1_N(_12017_),
    .X(_12192_));
 sky130_fd_sc_hd__xor2_2 _22520_ (.A(_12191_),
    .B(_12192_),
    .X(_12193_));
 sky130_fd_sc_hd__a21oi_2 _22521_ (.A1(_12023_),
    .A2(_12046_),
    .B1(_12193_),
    .Y(_12194_));
 sky130_fd_sc_hd__and3_2 _22522_ (.A(_12023_),
    .B(_12046_),
    .C(_12193_),
    .X(_12195_));
 sky130_fd_sc_hd__or2_2 _22523_ (.A(_12194_),
    .B(_12195_),
    .X(_12197_));
 sky130_fd_sc_hd__a31o_2 _22524_ (.A1(iX[4]),
    .A2(iY[31]),
    .A3(_11991_),
    .B1(_11989_),
    .X(_12198_));
 sky130_fd_sc_hd__xor2_2 _22525_ (.A(_12197_),
    .B(_12198_),
    .X(_12199_));
 sky130_fd_sc_hd__a21oi_2 _22526_ (.A1(_12028_),
    .A2(_12045_),
    .B1(_12199_),
    .Y(_12200_));
 sky130_fd_sc_hd__and3_2 _22527_ (.A(_12028_),
    .B(_12045_),
    .C(_12199_),
    .X(_12201_));
 sky130_fd_sc_hd__or2_2 _22528_ (.A(_12200_),
    .B(_12201_),
    .X(_12202_));
 sky130_fd_sc_hd__nand2_2 _22529_ (.A(_11775_),
    .B(_12036_),
    .Y(_12203_));
 sky130_fd_sc_hd__a2111o_2 _22530_ (.A1(_11188_),
    .A2(_11185_),
    .B1(_11367_),
    .C1(_11559_),
    .D1(_12203_),
    .X(_12204_));
 sky130_fd_sc_hd__nor2_2 _22531_ (.A(_11364_),
    .B(_11557_),
    .Y(_12205_));
 sky130_fd_sc_hd__nor2_2 _22532_ (.A(_11773_),
    .B(_12035_),
    .Y(_12206_));
 sky130_fd_sc_hd__nor2_2 _22533_ (.A(_12034_),
    .B(_12206_),
    .Y(_12208_));
 sky130_fd_sc_hd__o31a_2 _22534_ (.A1(_11558_),
    .A2(_12203_),
    .A3(_12205_),
    .B1(_12208_),
    .X(_12209_));
 sky130_fd_sc_hd__nand2_2 _22535_ (.A(_12204_),
    .B(_12209_),
    .Y(_12210_));
 sky130_fd_sc_hd__xnor2_2 _22536_ (.A(_12202_),
    .B(_12210_),
    .Y(_12211_));
 sky130_fd_sc_hd__nand2_2 _22537_ (.A(_11797_),
    .B(_11844_),
    .Y(_12212_));
 sky130_fd_sc_hd__and2b_2 _22538_ (.A_N(_11833_),
    .B(_11836_),
    .X(_12213_));
 sky130_fd_sc_hd__nor2_2 _22539_ (.A(_11837_),
    .B(_11843_),
    .Y(_12214_));
 sky130_fd_sc_hd__and2_2 _22540_ (.A(iX[4]),
    .B(iX[36]),
    .X(_12215_));
 sky130_fd_sc_hd__nor2_2 _22541_ (.A(iX[4]),
    .B(iX[36]),
    .Y(_12216_));
 sky130_fd_sc_hd__nor2_4 _22542_ (.A(_12215_),
    .B(_12216_),
    .Y(_12217_));
 sky130_fd_sc_hd__and2_2 _22543_ (.A(_11782_),
    .B(_11823_),
    .X(_12219_));
 sky130_fd_sc_hd__and2_2 _22544_ (.A(_11825_),
    .B(_11823_),
    .X(_12220_));
 sky130_fd_sc_hd__and2_2 _22545_ (.A(iX[3]),
    .B(iX[35]),
    .X(_12221_));
 sky130_fd_sc_hd__a211o_4 _22546_ (.A1(_11780_),
    .A2(_12219_),
    .B1(_12220_),
    .C1(_12221_),
    .X(_12222_));
 sky130_fd_sc_hd__xnor2_2 _22547_ (.A(_12217_),
    .B(_12222_),
    .Y(_12223_));
 sky130_fd_sc_hd__or4_2 _22548_ (.A(_11565_),
    .B(_11574_),
    .C(_11827_),
    .D(_12223_),
    .X(_12224_));
 sky130_fd_sc_hd__xor2_2 _22549_ (.A(_12217_),
    .B(_12222_),
    .X(_12225_));
 sky130_fd_sc_hd__a22o_2 _22550_ (.A1(_11582_),
    .A2(_11829_),
    .B1(_12225_),
    .B2(_11379_),
    .X(_12226_));
 sky130_fd_sc_hd__xnor2_2 _22551_ (.A(_11780_),
    .B(_11782_),
    .Y(_12227_));
 sky130_fd_sc_hd__nor2_2 _22552_ (.A(_12227_),
    .B(_11791_),
    .Y(_12228_));
 sky130_fd_sc_hd__nand3_2 _22553_ (.A(_12224_),
    .B(_12226_),
    .C(_12228_),
    .Y(_12230_));
 sky130_fd_sc_hd__a21o_2 _22554_ (.A1(_12224_),
    .A2(_12226_),
    .B1(_12228_),
    .X(_12231_));
 sky130_fd_sc_hd__a21o_2 _22555_ (.A1(_11830_),
    .A2(_11832_),
    .B1(_11828_),
    .X(_12232_));
 sky130_fd_sc_hd__nand3_2 _22556_ (.A(_12230_),
    .B(_12231_),
    .C(_12232_),
    .Y(_12233_));
 sky130_fd_sc_hd__a21o_2 _22557_ (.A1(_12230_),
    .A2(_12231_),
    .B1(_12232_),
    .X(_12234_));
 sky130_fd_sc_hd__nand2_2 _22558_ (.A(_12233_),
    .B(_12234_),
    .Y(_12235_));
 sky130_fd_sc_hd__and2_2 _22559_ (.A(iY[4]),
    .B(iY[36]),
    .X(_12236_));
 sky130_fd_sc_hd__nor2_2 _22560_ (.A(iY[4]),
    .B(iY[36]),
    .Y(_12237_));
 sky130_fd_sc_hd__nor2_2 _22561_ (.A(_12236_),
    .B(_12237_),
    .Y(_12238_));
 sky130_fd_sc_hd__a21boi_4 _22562_ (.A1(_11839_),
    .A2(_11841_),
    .B1_N(_11838_),
    .Y(_12239_));
 sky130_fd_sc_hd__xnor2_2 _22563_ (.A(_12238_),
    .B(_12239_),
    .Y(_12241_));
 sky130_fd_sc_hd__buf_1 _22564_ (.A(_12241_),
    .X(_12242_));
 sky130_fd_sc_hd__buf_1 _22565_ (.A(_12242_),
    .X(_12243_));
 sky130_fd_sc_hd__xor2_2 _22566_ (.A(_11840_),
    .B(_11841_),
    .X(_12244_));
 sky130_fd_sc_hd__nor2_2 _22567_ (.A(_11569_),
    .B(_12244_),
    .Y(_12245_));
 sky130_fd_sc_hd__a21o_2 _22568_ (.A1(_11374_),
    .A2(_12243_),
    .B1(_12245_),
    .X(_12246_));
 sky130_fd_sc_hd__xor2_2 _22569_ (.A(_12238_),
    .B(_12239_),
    .X(_12247_));
 sky130_fd_sc_hd__buf_1 _22570_ (.A(_12247_),
    .X(_12248_));
 sky130_fd_sc_hd__or3_2 _22571_ (.A(_11570_),
    .B(_11843_),
    .C(_12248_),
    .X(_12249_));
 sky130_fd_sc_hd__nand2_2 _22572_ (.A(_12246_),
    .B(_12249_),
    .Y(_12250_));
 sky130_fd_sc_hd__xor2_2 _22573_ (.A(_12235_),
    .B(_12250_),
    .X(_12252_));
 sky130_fd_sc_hd__o21a_2 _22574_ (.A1(_12213_),
    .A2(_12214_),
    .B1(_12252_),
    .X(_12253_));
 sky130_fd_sc_hd__nor3_2 _22575_ (.A(_12213_),
    .B(_12214_),
    .C(_12252_),
    .Y(_12254_));
 sky130_fd_sc_hd__or2_2 _22576_ (.A(_12253_),
    .B(_12254_),
    .X(_12255_));
 sky130_fd_sc_hd__xor2_2 _22577_ (.A(_12212_),
    .B(_12255_),
    .X(_12256_));
 sky130_fd_sc_hd__nand2_2 _22578_ (.A(_11801_),
    .B(_11851_),
    .Y(_12257_));
 sky130_fd_sc_hd__and3_2 _22579_ (.A(iX[33]),
    .B(iX[34]),
    .C(iY[35]),
    .X(_12258_));
 sky130_fd_sc_hd__a22o_2 _22580_ (.A1(iX[34]),
    .A2(iY[34]),
    .B1(iY[35]),
    .B2(iX[33]),
    .X(_12259_));
 sky130_fd_sc_hd__a21bo_2 _22581_ (.A1(iY[34]),
    .A2(_12258_),
    .B1_N(_12259_),
    .X(_12260_));
 sky130_fd_sc_hd__nand2_2 _22582_ (.A(iY[33]),
    .B(iX[35]),
    .Y(_12261_));
 sky130_fd_sc_hd__xor2_2 _22583_ (.A(_12260_),
    .B(_12261_),
    .X(_12263_));
 sky130_fd_sc_hd__a31o_2 _22584_ (.A1(iY[33]),
    .A2(iX[34]),
    .A3(_11848_),
    .B1(_11847_),
    .X(_12264_));
 sky130_fd_sc_hd__xor2_2 _22585_ (.A(_12263_),
    .B(_12264_),
    .X(_12265_));
 sky130_fd_sc_hd__a22oi_2 _22586_ (.A1(iY[32]),
    .A2(iX[36]),
    .B1(iY[36]),
    .B2(iX[32]),
    .Y(_12266_));
 sky130_fd_sc_hd__and4_2 _22587_ (.A(iX[32]),
    .B(iY[32]),
    .C(iX[36]),
    .D(iY[36]),
    .X(_12267_));
 sky130_fd_sc_hd__nor2_2 _22588_ (.A(_12266_),
    .B(_12267_),
    .Y(_12268_));
 sky130_fd_sc_hd__xnor2_2 _22589_ (.A(_12265_),
    .B(_12268_),
    .Y(_12269_));
 sky130_fd_sc_hd__a21oi_2 _22590_ (.A1(_12257_),
    .A2(_11854_),
    .B1(_12269_),
    .Y(_12270_));
 sky130_fd_sc_hd__and3_2 _22591_ (.A(_12257_),
    .B(_11854_),
    .C(_12269_),
    .X(_12271_));
 sky130_fd_sc_hd__nor2_2 _22592_ (.A(_12270_),
    .B(_12271_),
    .Y(_12272_));
 sky130_fd_sc_hd__or3_2 _22593_ (.A(_11856_),
    .B(_11861_),
    .C(_12272_),
    .X(_12274_));
 sky130_fd_sc_hd__nand2_2 _22594_ (.A(_11856_),
    .B(_12272_),
    .Y(_12275_));
 sky130_fd_sc_hd__nand2_2 _22595_ (.A(_11861_),
    .B(_12272_),
    .Y(_12276_));
 sky130_fd_sc_hd__and3_2 _22596_ (.A(_12274_),
    .B(_12275_),
    .C(_12276_),
    .X(_12277_));
 sky130_fd_sc_hd__xnor2_2 _22597_ (.A(_12256_),
    .B(_12277_),
    .Y(_12278_));
 sky130_fd_sc_hd__xnor2_2 _22598_ (.A(_11300_),
    .B(_12278_),
    .Y(_12279_));
 sky130_fd_sc_hd__or2_2 _22599_ (.A(_11845_),
    .B(_11863_),
    .X(_12280_));
 sky130_fd_sc_hd__o21a_2 _22600_ (.A1(oO[3]),
    .A2(_11864_),
    .B1(_12280_),
    .X(_12281_));
 sky130_fd_sc_hd__xnor2_2 _22601_ (.A(_12279_),
    .B(_12281_),
    .Y(_12282_));
 sky130_fd_sc_hd__a21o_2 _22602_ (.A1(_11865_),
    .A2(_11866_),
    .B1(_11870_),
    .X(_12283_));
 sky130_fd_sc_hd__xnor2_2 _22603_ (.A(_12282_),
    .B(_12283_),
    .Y(_12285_));
 sky130_fd_sc_hd__and2_2 _22604_ (.A(_12211_),
    .B(_12285_),
    .X(_12286_));
 sky130_fd_sc_hd__nor2_2 _22605_ (.A(_12211_),
    .B(_12285_),
    .Y(_12287_));
 sky130_fd_sc_hd__or2_2 _22606_ (.A(_12286_),
    .B(_12287_),
    .X(_12288_));
 sky130_fd_sc_hd__o21ba_2 _22607_ (.A1(_12041_),
    .A2(_12044_),
    .B1_N(_12040_),
    .X(_12289_));
 sky130_fd_sc_hd__nor2_2 _22608_ (.A(_12288_),
    .B(_12289_),
    .Y(_12290_));
 sky130_fd_sc_hd__and2_2 _22609_ (.A(_12288_),
    .B(_12289_),
    .X(_12291_));
 sky130_fd_sc_hd__nor2_2 _22610_ (.A(_12290_),
    .B(_12291_),
    .Y(oO[36]));
 sky130_fd_sc_hd__or2_2 _22611_ (.A(_12286_),
    .B(_12290_),
    .X(_12292_));
 sky130_fd_sc_hd__and2b_2 _22612_ (.A_N(_12197_),
    .B(_12198_),
    .X(_12293_));
 sky130_fd_sc_hd__nand2_2 _22613_ (.A(iY[7]),
    .B(iX[31]),
    .Y(_12295_));
 sky130_fd_sc_hd__and2_2 _22614_ (.A(iY[7]),
    .B(iX[30]),
    .X(_12296_));
 sky130_fd_sc_hd__a21o_2 _22615_ (.A1(iY[6]),
    .A2(iX[31]),
    .B1(_12296_),
    .X(_12297_));
 sky130_fd_sc_hd__o21ai_2 _22616_ (.A1(_12052_),
    .A2(_12295_),
    .B1(_12297_),
    .Y(_12298_));
 sky130_fd_sc_hd__nand2_2 _22617_ (.A(iY[8]),
    .B(iX[29]),
    .Y(_12299_));
 sky130_fd_sc_hd__xor2_2 _22618_ (.A(_12298_),
    .B(_12299_),
    .X(_12300_));
 sky130_fd_sc_hd__o21ai_2 _22619_ (.A1(_12051_),
    .A2(_12055_),
    .B1(_12300_),
    .Y(_12301_));
 sky130_fd_sc_hd__or3_2 _22620_ (.A(_12051_),
    .B(_12055_),
    .C(_12300_),
    .X(_12302_));
 sky130_fd_sc_hd__nand2_2 _22621_ (.A(_12301_),
    .B(_12302_),
    .Y(_12303_));
 sky130_fd_sc_hd__or2_2 _22622_ (.A(_12062_),
    .B(_12303_),
    .X(_12304_));
 sky130_fd_sc_hd__nand2_2 _22623_ (.A(_12062_),
    .B(_12303_),
    .Y(_12306_));
 sky130_fd_sc_hd__and2_2 _22624_ (.A(_12304_),
    .B(_12306_),
    .X(_12307_));
 sky130_fd_sc_hd__and2b_2 _22625_ (.A_N(_12080_),
    .B(_12079_),
    .X(_12308_));
 sky130_fd_sc_hd__or2b_2 _22626_ (.A(_12060_),
    .B_N(_12049_),
    .X(_12309_));
 sky130_fd_sc_hd__and4_2 _22627_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[24]),
    .D(iX[25]),
    .X(_12310_));
 sky130_fd_sc_hd__a22oi_2 _22628_ (.A1(iY[13]),
    .A2(iX[24]),
    .B1(iX[25]),
    .B2(iY[12]),
    .Y(_12311_));
 sky130_fd_sc_hd__nor2_2 _22629_ (.A(_12310_),
    .B(_12311_),
    .Y(_12312_));
 sky130_fd_sc_hd__nand2_2 _22630_ (.A(iY[14]),
    .B(iX[23]),
    .Y(_12313_));
 sky130_fd_sc_hd__xnor2_2 _22631_ (.A(_12312_),
    .B(_12313_),
    .Y(_12314_));
 sky130_fd_sc_hd__and4_2 _22632_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[27]),
    .D(iX[28]),
    .X(_12315_));
 sky130_fd_sc_hd__a22oi_2 _22633_ (.A1(iY[10]),
    .A2(iX[27]),
    .B1(iX[28]),
    .B2(iY[9]),
    .Y(_12317_));
 sky130_fd_sc_hd__nor2_2 _22634_ (.A(_12315_),
    .B(_12317_),
    .Y(_12318_));
 sky130_fd_sc_hd__nand2_2 _22635_ (.A(iY[11]),
    .B(iX[26]),
    .Y(_12319_));
 sky130_fd_sc_hd__xnor2_2 _22636_ (.A(_12318_),
    .B(_12319_),
    .Y(_12320_));
 sky130_fd_sc_hd__o21ba_2 _22637_ (.A1(_12076_),
    .A2(_12078_),
    .B1_N(_12074_),
    .X(_12321_));
 sky130_fd_sc_hd__xnor2_2 _22638_ (.A(_12320_),
    .B(_12321_),
    .Y(_12322_));
 sky130_fd_sc_hd__and2_2 _22639_ (.A(_12314_),
    .B(_12322_),
    .X(_12323_));
 sky130_fd_sc_hd__nor2_2 _22640_ (.A(_12314_),
    .B(_12322_),
    .Y(_12324_));
 sky130_fd_sc_hd__or2_2 _22641_ (.A(_12323_),
    .B(_12324_),
    .X(_12325_));
 sky130_fd_sc_hd__a21o_2 _22642_ (.A1(_12058_),
    .A2(_12309_),
    .B1(_12325_),
    .X(_12326_));
 sky130_fd_sc_hd__nand3_2 _22643_ (.A(_12058_),
    .B(_12309_),
    .C(_12325_),
    .Y(_12328_));
 sky130_fd_sc_hd__o211ai_2 _22644_ (.A1(_12308_),
    .A2(_12082_),
    .B1(_12326_),
    .C1(_12328_),
    .Y(_12329_));
 sky130_fd_sc_hd__a211o_2 _22645_ (.A1(_12326_),
    .A2(_12328_),
    .B1(_12308_),
    .C1(_12082_),
    .X(_12330_));
 sky130_fd_sc_hd__nand3_2 _22646_ (.A(_12307_),
    .B(_12329_),
    .C(_12330_),
    .Y(_12331_));
 sky130_fd_sc_hd__a21o_2 _22647_ (.A1(_12329_),
    .A2(_12330_),
    .B1(_12307_),
    .X(_12332_));
 sky130_fd_sc_hd__and2_2 _22648_ (.A(_12331_),
    .B(_12332_),
    .X(_12333_));
 sky130_fd_sc_hd__or2b_2 _22649_ (.A(_11894_),
    .B_N(_12065_),
    .X(_12334_));
 sky130_fd_sc_hd__nand2_2 _22650_ (.A(_12334_),
    .B(_12090_),
    .Y(_12335_));
 sky130_fd_sc_hd__xnor2_2 _22651_ (.A(_12333_),
    .B(_12335_),
    .Y(_12336_));
 sky130_fd_sc_hd__inv_2 _22652_ (.A(_12124_),
    .Y(_12337_));
 sky130_fd_sc_hd__and4_2 _22653_ (.A(iX[15]),
    .B(iX[16]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_12338_));
 sky130_fd_sc_hd__a22oi_2 _22654_ (.A1(iX[16]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[15]),
    .Y(_12339_));
 sky130_fd_sc_hd__nor2_2 _22655_ (.A(_12338_),
    .B(_12339_),
    .Y(_12340_));
 sky130_fd_sc_hd__nand2_2 _22656_ (.A(iX[14]),
    .B(iY[23]),
    .Y(_12341_));
 sky130_fd_sc_hd__xnor2_2 _22657_ (.A(_12340_),
    .B(_12341_),
    .Y(_12342_));
 sky130_fd_sc_hd__and4_2 _22658_ (.A(iX[18]),
    .B(iY[18]),
    .C(iX[19]),
    .D(iY[19]),
    .X(_12343_));
 sky130_fd_sc_hd__a22oi_2 _22659_ (.A1(iY[18]),
    .A2(iX[19]),
    .B1(iY[19]),
    .B2(iX[18]),
    .Y(_12344_));
 sky130_fd_sc_hd__nor2_2 _22660_ (.A(_12343_),
    .B(_12344_),
    .Y(_12345_));
 sky130_fd_sc_hd__nand2_2 _22661_ (.A(iX[17]),
    .B(iY[20]),
    .Y(_12346_));
 sky130_fd_sc_hd__xnor2_2 _22662_ (.A(_12345_),
    .B(_12346_),
    .Y(_12347_));
 sky130_fd_sc_hd__o21ba_2 _22663_ (.A1(_12102_),
    .A2(_12104_),
    .B1_N(_12101_),
    .X(_12349_));
 sky130_fd_sc_hd__xnor2_2 _22664_ (.A(_12347_),
    .B(_12349_),
    .Y(_12350_));
 sky130_fd_sc_hd__and2_2 _22665_ (.A(_12342_),
    .B(_12350_),
    .X(_12351_));
 sky130_fd_sc_hd__nor2_2 _22666_ (.A(_12342_),
    .B(_12350_),
    .Y(_12352_));
 sky130_fd_sc_hd__or2_2 _22667_ (.A(_12351_),
    .B(_12352_),
    .X(_12353_));
 sky130_fd_sc_hd__or3_2 _22668_ (.A(_12113_),
    .B(_12116_),
    .C(_12117_),
    .X(_12354_));
 sky130_fd_sc_hd__o21ba_2 _22669_ (.A1(_12070_),
    .A2(_12072_),
    .B1_N(_12069_),
    .X(_12355_));
 sky130_fd_sc_hd__nand4_2 _22670_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[21]),
    .D(iX[22]),
    .Y(_12356_));
 sky130_fd_sc_hd__a22o_2 _22671_ (.A1(iY[16]),
    .A2(iX[21]),
    .B1(iX[22]),
    .B2(iY[15]),
    .X(_12357_));
 sky130_fd_sc_hd__and2_2 _22672_ (.A(iY[17]),
    .B(iX[20]),
    .X(_12358_));
 sky130_fd_sc_hd__a21oi_2 _22673_ (.A1(_12356_),
    .A2(_12357_),
    .B1(_12358_),
    .Y(_12360_));
 sky130_fd_sc_hd__and3_2 _22674_ (.A(_12356_),
    .B(_12357_),
    .C(_12358_),
    .X(_12361_));
 sky130_fd_sc_hd__nor2_2 _22675_ (.A(_12360_),
    .B(_12361_),
    .Y(_12362_));
 sky130_fd_sc_hd__xnor2_2 _22676_ (.A(_12355_),
    .B(_12362_),
    .Y(_12363_));
 sky130_fd_sc_hd__o21ai_2 _22677_ (.A1(_12114_),
    .A2(_12116_),
    .B1(_12363_),
    .Y(_12364_));
 sky130_fd_sc_hd__or3_2 _22678_ (.A(_12114_),
    .B(_12116_),
    .C(_12363_),
    .X(_12365_));
 sky130_fd_sc_hd__nand2_2 _22679_ (.A(_12364_),
    .B(_12365_),
    .Y(_12366_));
 sky130_fd_sc_hd__a21oi_2 _22680_ (.A1(_12354_),
    .A2(_12121_),
    .B1(_12366_),
    .Y(_12367_));
 sky130_fd_sc_hd__and3_2 _22681_ (.A(_12354_),
    .B(_12121_),
    .C(_12366_),
    .X(_12368_));
 sky130_fd_sc_hd__or3_2 _22682_ (.A(_12353_),
    .B(_12367_),
    .C(_12368_),
    .X(_12369_));
 sky130_fd_sc_hd__o21ai_2 _22683_ (.A1(_12367_),
    .A2(_12368_),
    .B1(_12353_),
    .Y(_12371_));
 sky130_fd_sc_hd__nand2_2 _22684_ (.A(_12369_),
    .B(_12371_),
    .Y(_12372_));
 sky130_fd_sc_hd__a21oi_2 _22685_ (.A1(_12085_),
    .A2(_12088_),
    .B1(_12372_),
    .Y(_12373_));
 sky130_fd_sc_hd__and3_2 _22686_ (.A(_12085_),
    .B(_12088_),
    .C(_12372_),
    .X(_12374_));
 sky130_fd_sc_hd__a211oi_2 _22687_ (.A1(_12337_),
    .A2(_12126_),
    .B1(_12373_),
    .C1(_12374_),
    .Y(_12375_));
 sky130_fd_sc_hd__o211a_2 _22688_ (.A1(_12373_),
    .A2(_12374_),
    .B1(_12337_),
    .C1(_12126_),
    .X(_12376_));
 sky130_fd_sc_hd__or3_2 _22689_ (.A(_12336_),
    .B(_12375_),
    .C(_12376_),
    .X(_12377_));
 sky130_fd_sc_hd__o21ai_2 _22690_ (.A1(_12375_),
    .A2(_12376_),
    .B1(_12336_),
    .Y(_12378_));
 sky130_fd_sc_hd__o211a_2 _22691_ (.A1(_12092_),
    .A2(_12134_),
    .B1(_12377_),
    .C1(_12378_),
    .X(_12379_));
 sky130_fd_sc_hd__a211oi_2 _22692_ (.A1(_12377_),
    .A2(_12378_),
    .B1(_12092_),
    .C1(_12134_),
    .Y(_12380_));
 sky130_fd_sc_hd__inv_2 _22693_ (.A(_12179_),
    .Y(_12382_));
 sky130_fd_sc_hd__or2b_2 _22694_ (.A(_12149_),
    .B_N(_12148_),
    .X(_12383_));
 sky130_fd_sc_hd__and4_2 _22695_ (.A(iX[9]),
    .B(iX[10]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_12384_));
 sky130_fd_sc_hd__a22oi_2 _22696_ (.A1(iX[10]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[9]),
    .Y(_12385_));
 sky130_fd_sc_hd__nor2_2 _22697_ (.A(_12384_),
    .B(_12385_),
    .Y(_12386_));
 sky130_fd_sc_hd__nand2_2 _22698_ (.A(iX[8]),
    .B(iY[29]),
    .Y(_12387_));
 sky130_fd_sc_hd__xnor2_2 _22699_ (.A(_12386_),
    .B(_12387_),
    .Y(_12388_));
 sky130_fd_sc_hd__o21ba_2 _22700_ (.A1(_12145_),
    .A2(_12147_),
    .B1_N(_12144_),
    .X(_12389_));
 sky130_fd_sc_hd__xnor2_2 _22701_ (.A(_12388_),
    .B(_12389_),
    .Y(_12390_));
 sky130_fd_sc_hd__nand2_2 _22702_ (.A(iX[7]),
    .B(iY[30]),
    .Y(_12391_));
 sky130_fd_sc_hd__xor2_2 _22703_ (.A(_12390_),
    .B(_12391_),
    .X(_12393_));
 sky130_fd_sc_hd__a21oi_2 _22704_ (.A1(_12383_),
    .A2(_12151_),
    .B1(_12393_),
    .Y(_12394_));
 sky130_fd_sc_hd__and3_2 _22705_ (.A(_12383_),
    .B(_12151_),
    .C(_12393_),
    .X(_12395_));
 sky130_fd_sc_hd__nor2_2 _22706_ (.A(_12394_),
    .B(_12395_),
    .Y(_12396_));
 sky130_fd_sc_hd__nand2_2 _22707_ (.A(iX[6]),
    .B(iY[31]),
    .Y(_12397_));
 sky130_fd_sc_hd__xnor2_2 _22708_ (.A(_12396_),
    .B(_12397_),
    .Y(_12398_));
 sky130_fd_sc_hd__or2b_2 _22709_ (.A(_12165_),
    .B_N(_12170_),
    .X(_12399_));
 sky130_fd_sc_hd__or2b_2 _22710_ (.A(_12164_),
    .B_N(_12171_),
    .X(_12400_));
 sky130_fd_sc_hd__and2b_2 _22711_ (.A_N(_12106_),
    .B(_12105_),
    .X(_12401_));
 sky130_fd_sc_hd__o21ba_2 _22712_ (.A1(_12167_),
    .A2(_12169_),
    .B1_N(_12166_),
    .X(_12402_));
 sky130_fd_sc_hd__o21ba_2 _22713_ (.A1(_12096_),
    .A2(_12099_),
    .B1_N(_12095_),
    .X(_12404_));
 sky130_fd_sc_hd__and4_2 _22714_ (.A(iX[12]),
    .B(iX[13]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_12405_));
 sky130_fd_sc_hd__a22oi_2 _22715_ (.A1(iX[13]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[12]),
    .Y(_12406_));
 sky130_fd_sc_hd__nor2_2 _22716_ (.A(_12405_),
    .B(_12406_),
    .Y(_12407_));
 sky130_fd_sc_hd__nand2_2 _22717_ (.A(iX[11]),
    .B(iY[26]),
    .Y(_12408_));
 sky130_fd_sc_hd__xnor2_2 _22718_ (.A(_12407_),
    .B(_12408_),
    .Y(_12409_));
 sky130_fd_sc_hd__xnor2_2 _22719_ (.A(_12404_),
    .B(_12409_),
    .Y(_12410_));
 sky130_fd_sc_hd__xnor2_2 _22720_ (.A(_12402_),
    .B(_12410_),
    .Y(_12411_));
 sky130_fd_sc_hd__o21a_2 _22721_ (.A1(_12401_),
    .A2(_12109_),
    .B1(_12411_),
    .X(_12412_));
 sky130_fd_sc_hd__nor3_2 _22722_ (.A(_12401_),
    .B(_12109_),
    .C(_12411_),
    .Y(_12413_));
 sky130_fd_sc_hd__a211oi_2 _22723_ (.A1(_12399_),
    .A2(_12400_),
    .B1(_12412_),
    .C1(_12413_),
    .Y(_12415_));
 sky130_fd_sc_hd__o211a_2 _22724_ (.A1(_12412_),
    .A2(_12413_),
    .B1(_12399_),
    .C1(_12400_),
    .X(_12416_));
 sky130_fd_sc_hd__nor2_2 _22725_ (.A(_12173_),
    .B(_12176_),
    .Y(_12417_));
 sky130_fd_sc_hd__or3_2 _22726_ (.A(_12415_),
    .B(_12416_),
    .C(_12417_),
    .X(_12418_));
 sky130_fd_sc_hd__o21ai_2 _22727_ (.A1(_12415_),
    .A2(_12416_),
    .B1(_12417_),
    .Y(_12419_));
 sky130_fd_sc_hd__and3_2 _22728_ (.A(_12398_),
    .B(_12418_),
    .C(_12419_),
    .X(_12420_));
 sky130_fd_sc_hd__a21oi_2 _22729_ (.A1(_12418_),
    .A2(_12419_),
    .B1(_12398_),
    .Y(_12421_));
 sky130_fd_sc_hd__nor2_2 _22730_ (.A(_12420_),
    .B(_12421_),
    .Y(_12422_));
 sky130_fd_sc_hd__o21ai_2 _22731_ (.A1(_12129_),
    .A2(_12132_),
    .B1(_12422_),
    .Y(_12423_));
 sky130_fd_sc_hd__or3_2 _22732_ (.A(_12129_),
    .B(_12132_),
    .C(_12422_),
    .X(_12424_));
 sky130_fd_sc_hd__o211ai_2 _22733_ (.A1(_12382_),
    .A2(_12181_),
    .B1(_12423_),
    .C1(_12424_),
    .Y(_12426_));
 sky130_fd_sc_hd__a211o_2 _22734_ (.A1(_12423_),
    .A2(_12424_),
    .B1(_12382_),
    .C1(_12181_),
    .X(_12427_));
 sky130_fd_sc_hd__and4bb_2 _22735_ (.A_N(_12379_),
    .B_N(_12380_),
    .C(_12426_),
    .D(_12427_),
    .X(_12428_));
 sky130_fd_sc_hd__a2bb2o_2 _22736_ (.A1_N(_12379_),
    .A2_N(_12380_),
    .B1(_12426_),
    .B2(_12427_),
    .X(_12429_));
 sky130_fd_sc_hd__and2b_2 _22737_ (.A_N(_12428_),
    .B(_12429_),
    .X(_12430_));
 sky130_fd_sc_hd__a21oi_2 _22738_ (.A1(_12139_),
    .A2(_12188_),
    .B1(_12137_),
    .Y(_12431_));
 sky130_fd_sc_hd__xnor2_2 _22739_ (.A(_12430_),
    .B(_12431_),
    .Y(_12432_));
 sky130_fd_sc_hd__o21ba_2 _22740_ (.A1(_12142_),
    .A2(_12186_),
    .B1_N(_12184_),
    .X(_12433_));
 sky130_fd_sc_hd__xnor2_2 _22741_ (.A(_12432_),
    .B(_12433_),
    .Y(_12434_));
 sky130_fd_sc_hd__and2b_2 _22742_ (.A_N(_12191_),
    .B(_12192_),
    .X(_12435_));
 sky130_fd_sc_hd__o21bai_2 _22743_ (.A1(_12189_),
    .A2(_12190_),
    .B1_N(_12435_),
    .Y(_12437_));
 sky130_fd_sc_hd__xnor2_2 _22744_ (.A(_12434_),
    .B(_12437_),
    .Y(_12438_));
 sky130_fd_sc_hd__a31o_2 _22745_ (.A1(iX[5]),
    .A2(iY[31]),
    .A3(_12157_),
    .B1(_12155_),
    .X(_12439_));
 sky130_fd_sc_hd__xnor2_2 _22746_ (.A(_12438_),
    .B(_12439_),
    .Y(_12440_));
 sky130_fd_sc_hd__o21ai_2 _22747_ (.A1(_12194_),
    .A2(_12293_),
    .B1(_12440_),
    .Y(_12441_));
 sky130_fd_sc_hd__inv_2 _22748_ (.A(_12441_),
    .Y(_12442_));
 sky130_fd_sc_hd__nor3_2 _22749_ (.A(_12194_),
    .B(_12293_),
    .C(_12440_),
    .Y(_12443_));
 sky130_fd_sc_hd__nor2_2 _22750_ (.A(_12442_),
    .B(_12443_),
    .Y(_12444_));
 sky130_fd_sc_hd__inv_2 _22751_ (.A(_12202_),
    .Y(_12445_));
 sky130_fd_sc_hd__a21oi_2 _22752_ (.A1(_12445_),
    .A2(_12210_),
    .B1(_12200_),
    .Y(_12446_));
 sky130_fd_sc_hd__xnor2_2 _22753_ (.A(_12444_),
    .B(_12446_),
    .Y(_12448_));
 sky130_fd_sc_hd__or2_2 _22754_ (.A(_12212_),
    .B(_12255_),
    .X(_12449_));
 sky130_fd_sc_hd__xor2_2 _22755_ (.A(_11788_),
    .B(_11790_),
    .X(_12450_));
 sky130_fd_sc_hd__buf_1 _22756_ (.A(_12450_),
    .X(_12451_));
 sky130_fd_sc_hd__nand2_2 _22757_ (.A(iX[5]),
    .B(iX[37]),
    .Y(_12452_));
 sky130_fd_sc_hd__or2_2 _22758_ (.A(iX[5]),
    .B(iX[37]),
    .X(_12453_));
 sky130_fd_sc_hd__and2_2 _22759_ (.A(_12452_),
    .B(_12453_),
    .X(_12454_));
 sky130_fd_sc_hd__a21oi_2 _22760_ (.A1(_12217_),
    .A2(_12222_),
    .B1(_12215_),
    .Y(_12455_));
 sky130_fd_sc_hd__xor2_2 _22761_ (.A(_12454_),
    .B(_12455_),
    .X(_12456_));
 sky130_fd_sc_hd__buf_1 _22762_ (.A(_12456_),
    .X(_12457_));
 sky130_fd_sc_hd__or4_2 _22763_ (.A(_11565_),
    .B(_11574_),
    .C(_12223_),
    .D(_12457_),
    .X(_12459_));
 sky130_fd_sc_hd__xnor2_2 _22764_ (.A(_12454_),
    .B(_12455_),
    .Y(_12460_));
 sky130_fd_sc_hd__a22o_2 _22765_ (.A1(_11582_),
    .A2(_12225_),
    .B1(_12460_),
    .B2(_11379_),
    .X(_12461_));
 sky130_fd_sc_hd__nand4_2 _22766_ (.A(_12451_),
    .B(_11829_),
    .C(_12459_),
    .D(_12461_),
    .Y(_12462_));
 sky130_fd_sc_hd__a22o_2 _22767_ (.A1(_12450_),
    .A2(_11829_),
    .B1(_12459_),
    .B2(_12461_),
    .X(_12463_));
 sky130_fd_sc_hd__nand2_2 _22768_ (.A(_12224_),
    .B(_12230_),
    .Y(_12464_));
 sky130_fd_sc_hd__and3_2 _22769_ (.A(_12462_),
    .B(_12463_),
    .C(_12464_),
    .X(_12465_));
 sky130_fd_sc_hd__a21oi_2 _22770_ (.A1(_12462_),
    .A2(_12463_),
    .B1(_12464_),
    .Y(_12466_));
 sky130_fd_sc_hd__and3_2 _22771_ (.A(_11783_),
    .B(_12245_),
    .C(_12241_),
    .X(_12467_));
 sky130_fd_sc_hd__buf_1 _22772_ (.A(_12227_),
    .X(_12468_));
 sky130_fd_sc_hd__o22a_2 _22773_ (.A1(_12468_),
    .A2(_12244_),
    .B1(_12247_),
    .B2(_11569_),
    .X(_12470_));
 sky130_fd_sc_hd__nor2_2 _22774_ (.A(_12467_),
    .B(_12470_),
    .Y(_12471_));
 sky130_fd_sc_hd__nand2_2 _22775_ (.A(iY[5]),
    .B(iY[37]),
    .Y(_12472_));
 sky130_fd_sc_hd__or2_2 _22776_ (.A(iY[5]),
    .B(iY[37]),
    .X(_12473_));
 sky130_fd_sc_hd__nand2_2 _22777_ (.A(_12472_),
    .B(_12473_),
    .Y(_12474_));
 sky130_fd_sc_hd__nand2_2 _22778_ (.A(iY[4]),
    .B(iY[36]),
    .Y(_12475_));
 sky130_fd_sc_hd__o21a_2 _22779_ (.A1(_12237_),
    .A2(_12239_),
    .B1(_12475_),
    .X(_12476_));
 sky130_fd_sc_hd__xor2_2 _22780_ (.A(_12474_),
    .B(_12476_),
    .X(_12477_));
 sky130_fd_sc_hd__nand2_2 _22781_ (.A(_11373_),
    .B(_12477_),
    .Y(_12478_));
 sky130_fd_sc_hd__xnor2_2 _22782_ (.A(_12471_),
    .B(_12478_),
    .Y(_12479_));
 sky130_fd_sc_hd__or3b_2 _22783_ (.A(_12465_),
    .B(_12466_),
    .C_N(_12479_),
    .X(_12481_));
 sky130_fd_sc_hd__o21bai_2 _22784_ (.A1(_12465_),
    .A2(_12466_),
    .B1_N(_12479_),
    .Y(_12482_));
 sky130_fd_sc_hd__o21ai_2 _22785_ (.A1(_12235_),
    .A2(_12250_),
    .B1(_12233_),
    .Y(_12483_));
 sky130_fd_sc_hd__and3_2 _22786_ (.A(_12481_),
    .B(_12482_),
    .C(_12483_),
    .X(_12484_));
 sky130_fd_sc_hd__a21oi_2 _22787_ (.A1(_12481_),
    .A2(_12482_),
    .B1(_12483_),
    .Y(_12485_));
 sky130_fd_sc_hd__or3_2 _22788_ (.A(_12249_),
    .B(_12484_),
    .C(_12485_),
    .X(_12486_));
 sky130_fd_sc_hd__o21ai_2 _22789_ (.A1(_12484_),
    .A2(_12485_),
    .B1(_12249_),
    .Y(_12487_));
 sky130_fd_sc_hd__and3_2 _22790_ (.A(_12253_),
    .B(_12486_),
    .C(_12487_),
    .X(_12488_));
 sky130_fd_sc_hd__a21oi_2 _22791_ (.A1(_12486_),
    .A2(_12487_),
    .B1(_12253_),
    .Y(_12489_));
 sky130_fd_sc_hd__nor3_2 _22792_ (.A(_12449_),
    .B(_12488_),
    .C(_12489_),
    .Y(_12490_));
 sky130_fd_sc_hd__o21a_2 _22793_ (.A1(_12488_),
    .A2(_12489_),
    .B1(_12449_),
    .X(_12492_));
 sky130_fd_sc_hd__nand2_2 _22794_ (.A(_12263_),
    .B(_12264_),
    .Y(_12493_));
 sky130_fd_sc_hd__nand2_2 _22795_ (.A(_12265_),
    .B(_12268_),
    .Y(_12494_));
 sky130_fd_sc_hd__and4_2 _22796_ (.A(iX[34]),
    .B(iY[34]),
    .C(iX[35]),
    .D(iY[35]),
    .X(_12495_));
 sky130_fd_sc_hd__a22oi_2 _22797_ (.A1(iY[34]),
    .A2(iX[35]),
    .B1(iY[35]),
    .B2(iX[34]),
    .Y(_12496_));
 sky130_fd_sc_hd__nand2_2 _22798_ (.A(iY[33]),
    .B(iX[36]),
    .Y(_12497_));
 sky130_fd_sc_hd__or3_2 _22799_ (.A(_12495_),
    .B(_12496_),
    .C(_12497_),
    .X(_12498_));
 sky130_fd_sc_hd__o21ai_2 _22800_ (.A1(_12495_),
    .A2(_12496_),
    .B1(_12497_),
    .Y(_12499_));
 sky130_fd_sc_hd__a32o_2 _22801_ (.A1(iY[33]),
    .A2(iX[35]),
    .A3(_12259_),
    .B1(_12258_),
    .B2(iY[34]),
    .X(_12500_));
 sky130_fd_sc_hd__and3_2 _22802_ (.A(_12498_),
    .B(_12499_),
    .C(_12500_),
    .X(_12501_));
 sky130_fd_sc_hd__a21o_2 _22803_ (.A1(_12498_),
    .A2(_12499_),
    .B1(_12500_),
    .X(_12503_));
 sky130_fd_sc_hd__and2b_2 _22804_ (.A_N(_12501_),
    .B(_12503_),
    .X(_12504_));
 sky130_fd_sc_hd__and4_2 _22805_ (.A(iX[33]),
    .B(iY[32]),
    .C(iY[36]),
    .D(iX[37]),
    .X(_12505_));
 sky130_fd_sc_hd__a22oi_2 _22806_ (.A1(iX[33]),
    .A2(iY[36]),
    .B1(iX[37]),
    .B2(iY[32]),
    .Y(_12506_));
 sky130_fd_sc_hd__nor2_2 _22807_ (.A(_12505_),
    .B(_12506_),
    .Y(_12507_));
 sky130_fd_sc_hd__nand2_2 _22808_ (.A(iX[32]),
    .B(iY[37]),
    .Y(_12508_));
 sky130_fd_sc_hd__xnor2_2 _22809_ (.A(_12507_),
    .B(_12508_),
    .Y(_12509_));
 sky130_fd_sc_hd__xnor2_2 _22810_ (.A(_12504_),
    .B(_12509_),
    .Y(_12510_));
 sky130_fd_sc_hd__a21oi_2 _22811_ (.A1(_12493_),
    .A2(_12494_),
    .B1(_12510_),
    .Y(_12511_));
 sky130_fd_sc_hd__nand3_2 _22812_ (.A(_12493_),
    .B(_12494_),
    .C(_12510_),
    .Y(_12512_));
 sky130_fd_sc_hd__or2b_2 _22813_ (.A(_12511_),
    .B_N(_12512_),
    .X(_12514_));
 sky130_fd_sc_hd__xor2_2 _22814_ (.A(_12267_),
    .B(_12514_),
    .X(_12515_));
 sky130_fd_sc_hd__inv_2 _22815_ (.A(_12270_),
    .Y(_12516_));
 sky130_fd_sc_hd__and2_2 _22816_ (.A(_12516_),
    .B(_12275_),
    .X(_12517_));
 sky130_fd_sc_hd__xnor2_2 _22817_ (.A(_12515_),
    .B(_12517_),
    .Y(_12518_));
 sky130_fd_sc_hd__nor2_2 _22818_ (.A(_12276_),
    .B(_12518_),
    .Y(_12519_));
 sky130_fd_sc_hd__and2_2 _22819_ (.A(_12276_),
    .B(_12518_),
    .X(_12520_));
 sky130_fd_sc_hd__nor2_2 _22820_ (.A(_12519_),
    .B(_12520_),
    .Y(_12521_));
 sky130_fd_sc_hd__or3_2 _22821_ (.A(_12490_),
    .B(_12492_),
    .C(_12521_),
    .X(_12522_));
 sky130_fd_sc_hd__o21ai_2 _22822_ (.A1(_12490_),
    .A2(_12492_),
    .B1(_12521_),
    .Y(_12523_));
 sky130_fd_sc_hd__nand3b_2 _22823_ (.A_N(oO[5]),
    .B(_12522_),
    .C(_12523_),
    .Y(_12525_));
 sky130_fd_sc_hd__a21bo_2 _22824_ (.A1(_12522_),
    .A2(_12523_),
    .B1_N(oO[5]),
    .X(_12526_));
 sky130_fd_sc_hd__and2_2 _22825_ (.A(_12525_),
    .B(_12526_),
    .X(_12527_));
 sky130_fd_sc_hd__and2b_2 _22826_ (.A_N(_12277_),
    .B(_12256_),
    .X(_12528_));
 sky130_fd_sc_hd__a21o_2 _22827_ (.A1(_11300_),
    .A2(_12278_),
    .B1(_12528_),
    .X(_12529_));
 sky130_fd_sc_hd__xor2_2 _22828_ (.A(_12527_),
    .B(_12529_),
    .X(_12530_));
 sky130_fd_sc_hd__or2b_2 _22829_ (.A(_12282_),
    .B_N(_12283_),
    .X(_12531_));
 sky130_fd_sc_hd__o21ai_2 _22830_ (.A1(_12279_),
    .A2(_12281_),
    .B1(_12531_),
    .Y(_12532_));
 sky130_fd_sc_hd__xor2_2 _22831_ (.A(_12530_),
    .B(_12532_),
    .X(_12533_));
 sky130_fd_sc_hd__or2_2 _22832_ (.A(_12448_),
    .B(_12533_),
    .X(_12534_));
 sky130_fd_sc_hd__and2_2 _22833_ (.A(_12448_),
    .B(_12533_),
    .X(_12536_));
 sky130_fd_sc_hd__inv_2 _22834_ (.A(_12536_),
    .Y(_12537_));
 sky130_fd_sc_hd__nand2_2 _22835_ (.A(_12534_),
    .B(_12537_),
    .Y(_12538_));
 sky130_fd_sc_hd__xnor2_2 _22836_ (.A(_12292_),
    .B(_12538_),
    .Y(oO[37]));
 sky130_fd_sc_hd__nand2_2 _22837_ (.A(_12434_),
    .B(_12437_),
    .Y(_12539_));
 sky130_fd_sc_hd__or2b_2 _22838_ (.A(_12438_),
    .B_N(_12439_),
    .X(_12540_));
 sky130_fd_sc_hd__and2b_2 _22839_ (.A_N(_12431_),
    .B(_12430_),
    .X(_12541_));
 sky130_fd_sc_hd__and2b_2 _22840_ (.A_N(_12433_),
    .B(_12432_),
    .X(_12542_));
 sky130_fd_sc_hd__nand2_2 _22841_ (.A(_12333_),
    .B(_12335_),
    .Y(_12543_));
 sky130_fd_sc_hd__inv_2 _22842_ (.A(_12367_),
    .Y(_12544_));
 sky130_fd_sc_hd__and4_2 _22843_ (.A(iX[16]),
    .B(iX[17]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_12546_));
 sky130_fd_sc_hd__a22oi_2 _22844_ (.A1(iX[17]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[16]),
    .Y(_12547_));
 sky130_fd_sc_hd__nor2_2 _22845_ (.A(_12546_),
    .B(_12547_),
    .Y(_12548_));
 sky130_fd_sc_hd__nand2_2 _22846_ (.A(iX[15]),
    .B(iY[23]),
    .Y(_12549_));
 sky130_fd_sc_hd__xnor2_2 _22847_ (.A(_12548_),
    .B(_12549_),
    .Y(_12550_));
 sky130_fd_sc_hd__and4_2 _22848_ (.A(iY[18]),
    .B(iX[19]),
    .C(iY[19]),
    .D(iX[20]),
    .X(_12551_));
 sky130_fd_sc_hd__a22oi_2 _22849_ (.A1(iX[19]),
    .A2(iY[19]),
    .B1(iX[20]),
    .B2(iY[18]),
    .Y(_12552_));
 sky130_fd_sc_hd__nor2_2 _22850_ (.A(_12551_),
    .B(_12552_),
    .Y(_12553_));
 sky130_fd_sc_hd__nand2_2 _22851_ (.A(iX[18]),
    .B(iY[20]),
    .Y(_12554_));
 sky130_fd_sc_hd__xnor2_2 _22852_ (.A(_12553_),
    .B(_12554_),
    .Y(_12555_));
 sky130_fd_sc_hd__o21ba_2 _22853_ (.A1(_12344_),
    .A2(_12346_),
    .B1_N(_12343_),
    .X(_12557_));
 sky130_fd_sc_hd__xnor2_2 _22854_ (.A(_12555_),
    .B(_12557_),
    .Y(_12558_));
 sky130_fd_sc_hd__and2_2 _22855_ (.A(_12550_),
    .B(_12558_),
    .X(_12559_));
 sky130_fd_sc_hd__nor2_2 _22856_ (.A(_12550_),
    .B(_12558_),
    .Y(_12560_));
 sky130_fd_sc_hd__or2_2 _22857_ (.A(_12559_),
    .B(_12560_),
    .X(_12561_));
 sky130_fd_sc_hd__or3_2 _22858_ (.A(_12355_),
    .B(_12360_),
    .C(_12361_),
    .X(_12562_));
 sky130_fd_sc_hd__and4_2 _22859_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[21]),
    .D(iX[22]),
    .X(_12563_));
 sky130_fd_sc_hd__o21ba_2 _22860_ (.A1(_12311_),
    .A2(_12313_),
    .B1_N(_12310_),
    .X(_12564_));
 sky130_fd_sc_hd__and4_2 _22861_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[22]),
    .D(iX[23]),
    .X(_12565_));
 sky130_fd_sc_hd__a22oi_2 _22862_ (.A1(iY[16]),
    .A2(iX[22]),
    .B1(iX[23]),
    .B2(iY[15]),
    .Y(_12566_));
 sky130_fd_sc_hd__nand2_2 _22863_ (.A(iY[17]),
    .B(iX[21]),
    .Y(_12568_));
 sky130_fd_sc_hd__o21a_2 _22864_ (.A1(_12565_),
    .A2(_12566_),
    .B1(_12568_),
    .X(_12569_));
 sky130_fd_sc_hd__nor3_2 _22865_ (.A(_12565_),
    .B(_12566_),
    .C(_12568_),
    .Y(_12570_));
 sky130_fd_sc_hd__nor2_2 _22866_ (.A(_12569_),
    .B(_12570_),
    .Y(_12571_));
 sky130_fd_sc_hd__xnor2_2 _22867_ (.A(_12564_),
    .B(_12571_),
    .Y(_12572_));
 sky130_fd_sc_hd__o21ai_2 _22868_ (.A1(_12563_),
    .A2(_12361_),
    .B1(_12572_),
    .Y(_12573_));
 sky130_fd_sc_hd__or3_2 _22869_ (.A(_12563_),
    .B(_12361_),
    .C(_12572_),
    .X(_12574_));
 sky130_fd_sc_hd__nand2_2 _22870_ (.A(_12573_),
    .B(_12574_),
    .Y(_12575_));
 sky130_fd_sc_hd__a21oi_2 _22871_ (.A1(_12562_),
    .A2(_12364_),
    .B1(_12575_),
    .Y(_12576_));
 sky130_fd_sc_hd__and3_2 _22872_ (.A(_12562_),
    .B(_12364_),
    .C(_12575_),
    .X(_12577_));
 sky130_fd_sc_hd__or3_2 _22873_ (.A(_12561_),
    .B(_12576_),
    .C(_12577_),
    .X(_12579_));
 sky130_fd_sc_hd__o21ai_2 _22874_ (.A1(_12576_),
    .A2(_12577_),
    .B1(_12561_),
    .Y(_12580_));
 sky130_fd_sc_hd__nand2_2 _22875_ (.A(_12579_),
    .B(_12580_),
    .Y(_12581_));
 sky130_fd_sc_hd__a21oi_2 _22876_ (.A1(_12326_),
    .A2(_12329_),
    .B1(_12581_),
    .Y(_12582_));
 sky130_fd_sc_hd__and3_2 _22877_ (.A(_12326_),
    .B(_12329_),
    .C(_12581_),
    .X(_12583_));
 sky130_fd_sc_hd__a211oi_2 _22878_ (.A1(_12544_),
    .A2(_12369_),
    .B1(_12582_),
    .C1(_12583_),
    .Y(_12584_));
 sky130_fd_sc_hd__o211a_2 _22879_ (.A1(_12582_),
    .A2(_12583_),
    .B1(_12544_),
    .C1(_12369_),
    .X(_12585_));
 sky130_fd_sc_hd__nand2_2 _22880_ (.A(iY[8]),
    .B(iX[31]),
    .Y(_12586_));
 sky130_fd_sc_hd__a22o_2 _22881_ (.A1(iY[8]),
    .A2(iX[30]),
    .B1(iX[31]),
    .B2(iY[7]),
    .X(_12587_));
 sky130_fd_sc_hd__o21a_2 _22882_ (.A1(_12050_),
    .A2(_12586_),
    .B1(_12587_),
    .X(_12588_));
 sky130_fd_sc_hd__o22ai_2 _22883_ (.A1(_12052_),
    .A2(_12295_),
    .B1(_12298_),
    .B2(_12299_),
    .Y(_12590_));
 sky130_fd_sc_hd__nand2_2 _22884_ (.A(_12588_),
    .B(_12590_),
    .Y(_12591_));
 sky130_fd_sc_hd__or2_2 _22885_ (.A(_12588_),
    .B(_12590_),
    .X(_12592_));
 sky130_fd_sc_hd__and2_2 _22886_ (.A(_12591_),
    .B(_12592_),
    .X(_12593_));
 sky130_fd_sc_hd__and2b_2 _22887_ (.A_N(_12321_),
    .B(_12320_),
    .X(_12594_));
 sky130_fd_sc_hd__and4_2 _22888_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[25]),
    .D(iX[26]),
    .X(_12595_));
 sky130_fd_sc_hd__a22oi_2 _22889_ (.A1(iY[13]),
    .A2(iX[25]),
    .B1(iX[26]),
    .B2(iY[12]),
    .Y(_12596_));
 sky130_fd_sc_hd__nor2_2 _22890_ (.A(_12595_),
    .B(_12596_),
    .Y(_12597_));
 sky130_fd_sc_hd__nand2_2 _22891_ (.A(iY[14]),
    .B(iX[24]),
    .Y(_12598_));
 sky130_fd_sc_hd__xnor2_2 _22892_ (.A(_12597_),
    .B(_12598_),
    .Y(_12599_));
 sky130_fd_sc_hd__and4_2 _22893_ (.A(iY[9]),
    .B(iY[10]),
    .C(iX[28]),
    .D(iX[29]),
    .X(_12601_));
 sky130_fd_sc_hd__and2_2 _22894_ (.A(iY[9]),
    .B(iX[29]),
    .X(_12602_));
 sky130_fd_sc_hd__a21oi_2 _22895_ (.A1(iY[10]),
    .A2(iX[28]),
    .B1(_12602_),
    .Y(_12603_));
 sky130_fd_sc_hd__nor2_2 _22896_ (.A(_12601_),
    .B(_12603_),
    .Y(_12604_));
 sky130_fd_sc_hd__nand2_2 _22897_ (.A(iY[11]),
    .B(iX[27]),
    .Y(_12605_));
 sky130_fd_sc_hd__xnor2_2 _22898_ (.A(_12604_),
    .B(_12605_),
    .Y(_12606_));
 sky130_fd_sc_hd__o21ba_2 _22899_ (.A1(_12317_),
    .A2(_12319_),
    .B1_N(_12315_),
    .X(_12607_));
 sky130_fd_sc_hd__xnor2_2 _22900_ (.A(_12606_),
    .B(_12607_),
    .Y(_12608_));
 sky130_fd_sc_hd__xnor2_2 _22901_ (.A(_12599_),
    .B(_12608_),
    .Y(_12609_));
 sky130_fd_sc_hd__or2_2 _22902_ (.A(_12301_),
    .B(_12609_),
    .X(_12610_));
 sky130_fd_sc_hd__nand2_2 _22903_ (.A(_12301_),
    .B(_12609_),
    .Y(_12612_));
 sky130_fd_sc_hd__and2_2 _22904_ (.A(_12610_),
    .B(_12612_),
    .X(_12613_));
 sky130_fd_sc_hd__o21ai_2 _22905_ (.A1(_12594_),
    .A2(_12323_),
    .B1(_12613_),
    .Y(_12614_));
 sky130_fd_sc_hd__or3_2 _22906_ (.A(_12594_),
    .B(_12323_),
    .C(_12613_),
    .X(_12615_));
 sky130_fd_sc_hd__and3_2 _22907_ (.A(_12593_),
    .B(_12614_),
    .C(_12615_),
    .X(_12616_));
 sky130_fd_sc_hd__a21oi_2 _22908_ (.A1(_12614_),
    .A2(_12615_),
    .B1(_12593_),
    .Y(_12617_));
 sky130_fd_sc_hd__a211o_2 _22909_ (.A1(_12304_),
    .A2(_12331_),
    .B1(_12616_),
    .C1(_12617_),
    .X(_12618_));
 sky130_fd_sc_hd__o211ai_2 _22910_ (.A1(_12616_),
    .A2(_12617_),
    .B1(_12304_),
    .C1(_12331_),
    .Y(_12619_));
 sky130_fd_sc_hd__nand2_2 _22911_ (.A(_12618_),
    .B(_12619_),
    .Y(_12620_));
 sky130_fd_sc_hd__o21a_2 _22912_ (.A1(_12584_),
    .A2(_12585_),
    .B1(_12620_),
    .X(_12621_));
 sky130_fd_sc_hd__or3_2 _22913_ (.A(_12620_),
    .B(_12584_),
    .C(_12585_),
    .X(_12623_));
 sky130_fd_sc_hd__inv_2 _22914_ (.A(_12623_),
    .Y(_12624_));
 sky130_fd_sc_hd__a211o_2 _22915_ (.A1(_12543_),
    .A2(_12377_),
    .B1(_12621_),
    .C1(_12624_),
    .X(_12625_));
 sky130_fd_sc_hd__o211ai_2 _22916_ (.A1(_12621_),
    .A2(_12624_),
    .B1(_12543_),
    .C1(_12377_),
    .Y(_12626_));
 sky130_fd_sc_hd__inv_2 _22917_ (.A(_12418_),
    .Y(_12627_));
 sky130_fd_sc_hd__and4_2 _22918_ (.A(iX[10]),
    .B(iX[11]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_12628_));
 sky130_fd_sc_hd__a22oi_2 _22919_ (.A1(iX[11]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[10]),
    .Y(_12629_));
 sky130_fd_sc_hd__nor2_2 _22920_ (.A(_12628_),
    .B(_12629_),
    .Y(_12630_));
 sky130_fd_sc_hd__nand2_2 _22921_ (.A(iX[9]),
    .B(iY[29]),
    .Y(_12631_));
 sky130_fd_sc_hd__xnor2_2 _22922_ (.A(_12630_),
    .B(_12631_),
    .Y(_12632_));
 sky130_fd_sc_hd__o21ba_2 _22923_ (.A1(_12385_),
    .A2(_12387_),
    .B1_N(_12384_),
    .X(_12634_));
 sky130_fd_sc_hd__xnor2_2 _22924_ (.A(_12632_),
    .B(_12634_),
    .Y(_12635_));
 sky130_fd_sc_hd__and2_2 _22925_ (.A(iX[8]),
    .B(iY[30]),
    .X(_12636_));
 sky130_fd_sc_hd__or2_2 _22926_ (.A(_12635_),
    .B(_12636_),
    .X(_12637_));
 sky130_fd_sc_hd__nand2_2 _22927_ (.A(_12635_),
    .B(_12636_),
    .Y(_12638_));
 sky130_fd_sc_hd__and2b_2 _22928_ (.A_N(_12389_),
    .B(_12388_),
    .X(_12639_));
 sky130_fd_sc_hd__a31o_2 _22929_ (.A1(iX[7]),
    .A2(iY[30]),
    .A3(_12390_),
    .B1(_12639_),
    .X(_12640_));
 sky130_fd_sc_hd__nand3_2 _22930_ (.A(_12637_),
    .B(_12638_),
    .C(_12640_),
    .Y(_12641_));
 sky130_fd_sc_hd__a21o_2 _22931_ (.A1(_12637_),
    .A2(_12638_),
    .B1(_12640_),
    .X(_12642_));
 sky130_fd_sc_hd__nand2_2 _22932_ (.A(_12641_),
    .B(_12642_),
    .Y(_12643_));
 sky130_fd_sc_hd__nand2_2 _22933_ (.A(iX[7]),
    .B(iY[31]),
    .Y(_12645_));
 sky130_fd_sc_hd__nand2_2 _22934_ (.A(_12643_),
    .B(_12645_),
    .Y(_12646_));
 sky130_fd_sc_hd__or2_2 _22935_ (.A(_12643_),
    .B(_12645_),
    .X(_12647_));
 sky130_fd_sc_hd__and2_2 _22936_ (.A(_12646_),
    .B(_12647_),
    .X(_12648_));
 sky130_fd_sc_hd__or2b_2 _22937_ (.A(_12404_),
    .B_N(_12409_),
    .X(_12649_));
 sky130_fd_sc_hd__or2b_2 _22938_ (.A(_12402_),
    .B_N(_12410_),
    .X(_12650_));
 sky130_fd_sc_hd__and2b_2 _22939_ (.A_N(_12349_),
    .B(_12347_),
    .X(_12651_));
 sky130_fd_sc_hd__o21ba_2 _22940_ (.A1(_12406_),
    .A2(_12408_),
    .B1_N(_12405_),
    .X(_12652_));
 sky130_fd_sc_hd__o21ba_2 _22941_ (.A1(_12339_),
    .A2(_12341_),
    .B1_N(_12338_),
    .X(_12653_));
 sky130_fd_sc_hd__and4_2 _22942_ (.A(iX[13]),
    .B(iX[14]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_12654_));
 sky130_fd_sc_hd__a22oi_2 _22943_ (.A1(iX[14]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[13]),
    .Y(_12656_));
 sky130_fd_sc_hd__nor2_2 _22944_ (.A(_12654_),
    .B(_12656_),
    .Y(_12657_));
 sky130_fd_sc_hd__nand2_2 _22945_ (.A(iX[12]),
    .B(iY[26]),
    .Y(_12658_));
 sky130_fd_sc_hd__xnor2_2 _22946_ (.A(_12657_),
    .B(_12658_),
    .Y(_12659_));
 sky130_fd_sc_hd__xnor2_2 _22947_ (.A(_12653_),
    .B(_12659_),
    .Y(_12660_));
 sky130_fd_sc_hd__xnor2_2 _22948_ (.A(_12652_),
    .B(_12660_),
    .Y(_12661_));
 sky130_fd_sc_hd__o21a_2 _22949_ (.A1(_12651_),
    .A2(_12351_),
    .B1(_12661_),
    .X(_12662_));
 sky130_fd_sc_hd__nor3_2 _22950_ (.A(_12651_),
    .B(_12351_),
    .C(_12661_),
    .Y(_12663_));
 sky130_fd_sc_hd__a211oi_2 _22951_ (.A1(_12649_),
    .A2(_12650_),
    .B1(_12662_),
    .C1(_12663_),
    .Y(_12664_));
 sky130_fd_sc_hd__o211a_2 _22952_ (.A1(_12662_),
    .A2(_12663_),
    .B1(_12649_),
    .C1(_12650_),
    .X(_12665_));
 sky130_fd_sc_hd__nor2_2 _22953_ (.A(_12412_),
    .B(_12415_),
    .Y(_12667_));
 sky130_fd_sc_hd__or3_2 _22954_ (.A(_12664_),
    .B(_12665_),
    .C(_12667_),
    .X(_12668_));
 sky130_fd_sc_hd__o21ai_2 _22955_ (.A1(_12664_),
    .A2(_12665_),
    .B1(_12667_),
    .Y(_12669_));
 sky130_fd_sc_hd__and3_2 _22956_ (.A(_12648_),
    .B(_12668_),
    .C(_12669_),
    .X(_12670_));
 sky130_fd_sc_hd__a21oi_2 _22957_ (.A1(_12668_),
    .A2(_12669_),
    .B1(_12648_),
    .Y(_12671_));
 sky130_fd_sc_hd__nor2_2 _22958_ (.A(_12670_),
    .B(_12671_),
    .Y(_12672_));
 sky130_fd_sc_hd__o21ai_2 _22959_ (.A1(_12373_),
    .A2(_12375_),
    .B1(_12672_),
    .Y(_12673_));
 sky130_fd_sc_hd__or3_2 _22960_ (.A(_12373_),
    .B(_12375_),
    .C(_12672_),
    .X(_12674_));
 sky130_fd_sc_hd__o211ai_2 _22961_ (.A1(_12627_),
    .A2(_12420_),
    .B1(_12673_),
    .C1(_12674_),
    .Y(_12675_));
 sky130_fd_sc_hd__a211o_2 _22962_ (.A1(_12673_),
    .A2(_12674_),
    .B1(_12627_),
    .C1(_12420_),
    .X(_12676_));
 sky130_fd_sc_hd__nand4_2 _22963_ (.A(_12625_),
    .B(_12626_),
    .C(_12675_),
    .D(_12676_),
    .Y(_12678_));
 sky130_fd_sc_hd__a22o_2 _22964_ (.A1(_12625_),
    .A2(_12626_),
    .B1(_12675_),
    .B2(_12676_),
    .X(_12679_));
 sky130_fd_sc_hd__o211a_2 _22965_ (.A1(_12379_),
    .A2(_12428_),
    .B1(_12678_),
    .C1(_12679_),
    .X(_12680_));
 sky130_fd_sc_hd__a211oi_2 _22966_ (.A1(_12678_),
    .A2(_12679_),
    .B1(_12379_),
    .C1(_12428_),
    .Y(_12681_));
 sky130_fd_sc_hd__or2_2 _22967_ (.A(_12680_),
    .B(_12681_),
    .X(_12682_));
 sky130_fd_sc_hd__nand2_2 _22968_ (.A(_12423_),
    .B(_12426_),
    .Y(_12683_));
 sky130_fd_sc_hd__xnor2_2 _22969_ (.A(_12682_),
    .B(_12683_),
    .Y(_12684_));
 sky130_fd_sc_hd__o21ai_2 _22970_ (.A1(_12541_),
    .A2(_12542_),
    .B1(_12684_),
    .Y(_12685_));
 sky130_fd_sc_hd__or3_2 _22971_ (.A(_12541_),
    .B(_12542_),
    .C(_12684_),
    .X(_12686_));
 sky130_fd_sc_hd__nand2_2 _22972_ (.A(_12685_),
    .B(_12686_),
    .Y(_12687_));
 sky130_fd_sc_hd__a31o_2 _22973_ (.A1(iX[6]),
    .A2(iY[31]),
    .A3(_12396_),
    .B1(_12394_),
    .X(_12689_));
 sky130_fd_sc_hd__xor2_2 _22974_ (.A(_12687_),
    .B(_12689_),
    .X(_12690_));
 sky130_fd_sc_hd__a21oi_2 _22975_ (.A1(_12539_),
    .A2(_12540_),
    .B1(_12690_),
    .Y(_12691_));
 sky130_fd_sc_hd__and3_2 _22976_ (.A(_12539_),
    .B(_12540_),
    .C(_12690_),
    .X(_12692_));
 sky130_fd_sc_hd__or2_2 _22977_ (.A(_12691_),
    .B(_12692_),
    .X(_12693_));
 sky130_fd_sc_hd__o21ai_2 _22978_ (.A1(_12443_),
    .A2(_12446_),
    .B1(_12441_),
    .Y(_12694_));
 sky130_fd_sc_hd__xnor2_2 _22979_ (.A(_12693_),
    .B(_12694_),
    .Y(_12695_));
 sky130_fd_sc_hd__nand2_2 _22980_ (.A(_12527_),
    .B(_12529_),
    .Y(_12696_));
 sky130_fd_sc_hd__nand2_2 _22981_ (.A(_12530_),
    .B(_12532_),
    .Y(_12697_));
 sky130_fd_sc_hd__and3b_2 _22982_ (.A_N(_12511_),
    .B(_12512_),
    .C(_12267_),
    .X(_12698_));
 sky130_fd_sc_hd__and4_2 _22983_ (.A(iY[34]),
    .B(iX[35]),
    .C(iY[35]),
    .D(iX[36]),
    .X(_12700_));
 sky130_fd_sc_hd__a22oi_2 _22984_ (.A1(iX[35]),
    .A2(iY[35]),
    .B1(iX[36]),
    .B2(iY[34]),
    .Y(_12701_));
 sky130_fd_sc_hd__nand2_2 _22985_ (.A(iY[33]),
    .B(iX[37]),
    .Y(_12702_));
 sky130_fd_sc_hd__or3_2 _22986_ (.A(_12700_),
    .B(_12701_),
    .C(_12702_),
    .X(_12703_));
 sky130_fd_sc_hd__o21ai_2 _22987_ (.A1(_12700_),
    .A2(_12701_),
    .B1(_12702_),
    .Y(_12704_));
 sky130_fd_sc_hd__o21bai_2 _22988_ (.A1(_12496_),
    .A2(_12497_),
    .B1_N(_12495_),
    .Y(_12705_));
 sky130_fd_sc_hd__nand3_2 _22989_ (.A(_12703_),
    .B(_12704_),
    .C(_12705_),
    .Y(_12706_));
 sky130_fd_sc_hd__a21o_2 _22990_ (.A1(_12703_),
    .A2(_12704_),
    .B1(_12705_),
    .X(_12707_));
 sky130_fd_sc_hd__and3_2 _22991_ (.A(iY[32]),
    .B(iX[34]),
    .C(iX[38]),
    .X(_12708_));
 sky130_fd_sc_hd__a22o_2 _22992_ (.A1(iX[34]),
    .A2(iY[36]),
    .B1(iX[38]),
    .B2(iY[32]),
    .X(_12709_));
 sky130_fd_sc_hd__a21bo_2 _22993_ (.A1(iY[36]),
    .A2(_12708_),
    .B1_N(_12709_),
    .X(_12711_));
 sky130_fd_sc_hd__nand2_2 _22994_ (.A(iX[33]),
    .B(iY[37]),
    .Y(_12712_));
 sky130_fd_sc_hd__xor2_2 _22995_ (.A(_12711_),
    .B(_12712_),
    .X(_12713_));
 sky130_fd_sc_hd__nand3_2 _22996_ (.A(_12706_),
    .B(_12707_),
    .C(_12713_),
    .Y(_12714_));
 sky130_fd_sc_hd__a21o_2 _22997_ (.A1(_12706_),
    .A2(_12707_),
    .B1(_12713_),
    .X(_12715_));
 sky130_fd_sc_hd__a21o_2 _22998_ (.A1(_12503_),
    .A2(_12509_),
    .B1(_12501_),
    .X(_12716_));
 sky130_fd_sc_hd__and3_2 _22999_ (.A(_12714_),
    .B(_12715_),
    .C(_12716_),
    .X(_12717_));
 sky130_fd_sc_hd__inv_2 _23000_ (.A(_12717_),
    .Y(_12718_));
 sky130_fd_sc_hd__a21o_2 _23001_ (.A1(_12714_),
    .A2(_12715_),
    .B1(_12716_),
    .X(_12719_));
 sky130_fd_sc_hd__and3_2 _23002_ (.A(iX[32]),
    .B(iY[37]),
    .C(_12507_),
    .X(_12720_));
 sky130_fd_sc_hd__o211a_2 _23003_ (.A1(_12505_),
    .A2(_12720_),
    .B1(iX[32]),
    .C1(iY[38]),
    .X(_12722_));
 sky130_fd_sc_hd__a211oi_2 _23004_ (.A1(iX[32]),
    .A2(iY[38]),
    .B1(_12505_),
    .C1(_12720_),
    .Y(_12723_));
 sky130_fd_sc_hd__nor2_2 _23005_ (.A(_12722_),
    .B(_12723_),
    .Y(_12724_));
 sky130_fd_sc_hd__nand3_2 _23006_ (.A(_12718_),
    .B(_12719_),
    .C(_12724_),
    .Y(_12725_));
 sky130_fd_sc_hd__a21o_2 _23007_ (.A1(_12718_),
    .A2(_12719_),
    .B1(_12724_),
    .X(_12726_));
 sky130_fd_sc_hd__o211ai_2 _23008_ (.A1(_12511_),
    .A2(_12698_),
    .B1(_12725_),
    .C1(_12726_),
    .Y(_12727_));
 sky130_fd_sc_hd__a211o_2 _23009_ (.A1(_12725_),
    .A2(_12726_),
    .B1(_12511_),
    .C1(_12698_),
    .X(_12728_));
 sky130_fd_sc_hd__and4bb_2 _23010_ (.A_N(_12516_),
    .B_N(_12515_),
    .C(_12727_),
    .D(_12728_),
    .X(_12729_));
 sky130_fd_sc_hd__o2bb2a_2 _23011_ (.A1_N(_12727_),
    .A2_N(_12728_),
    .B1(_12516_),
    .B2(_12515_),
    .X(_12730_));
 sky130_fd_sc_hd__nor2_2 _23012_ (.A(_12275_),
    .B(_12515_),
    .Y(_12731_));
 sky130_fd_sc_hd__or3b_2 _23013_ (.A(_12729_),
    .B(_12730_),
    .C_N(_12731_),
    .X(_12733_));
 sky130_fd_sc_hd__o21bai_2 _23014_ (.A1(_12729_),
    .A2(_12730_),
    .B1_N(_12731_),
    .Y(_12734_));
 sky130_fd_sc_hd__nand2_2 _23015_ (.A(_12733_),
    .B(_12734_),
    .Y(_12735_));
 sky130_fd_sc_hd__nor3_2 _23016_ (.A(_12276_),
    .B(_12518_),
    .C(_12735_),
    .Y(_12736_));
 sky130_fd_sc_hd__and2b_2 _23017_ (.A_N(_12519_),
    .B(_12735_),
    .X(_12737_));
 sky130_fd_sc_hd__nor2_2 _23018_ (.A(_12736_),
    .B(_12737_),
    .Y(_12738_));
 sky130_fd_sc_hd__nor2_2 _23019_ (.A(_11574_),
    .B(_12457_),
    .Y(_12739_));
 sky130_fd_sc_hd__and2_2 _23020_ (.A(iX[6]),
    .B(iX[38]),
    .X(_12740_));
 sky130_fd_sc_hd__nor2_2 _23021_ (.A(iX[6]),
    .B(iX[38]),
    .Y(_12741_));
 sky130_fd_sc_hd__nor2_2 _23022_ (.A(_12740_),
    .B(_12741_),
    .Y(_12742_));
 sky130_fd_sc_hd__or2b_2 _23023_ (.A(_12215_),
    .B_N(_12452_),
    .X(_12744_));
 sky130_fd_sc_hd__a21o_2 _23024_ (.A1(_12217_),
    .A2(_12222_),
    .B1(_12744_),
    .X(_12745_));
 sky130_fd_sc_hd__and3_2 _23025_ (.A(_12453_),
    .B(_12742_),
    .C(_12745_),
    .X(_12746_));
 sky130_fd_sc_hd__a21oi_2 _23026_ (.A1(_12453_),
    .A2(_12745_),
    .B1(_12742_),
    .Y(_12747_));
 sky130_fd_sc_hd__or3_2 _23027_ (.A(_11564_),
    .B(_12746_),
    .C(_12747_),
    .X(_12748_));
 sky130_fd_sc_hd__xnor2_2 _23028_ (.A(_12739_),
    .B(_12748_),
    .Y(_12749_));
 sky130_fd_sc_hd__nor2_2 _23029_ (.A(_11791_),
    .B(_12223_),
    .Y(_12750_));
 sky130_fd_sc_hd__xnor2_2 _23030_ (.A(_12749_),
    .B(_12750_),
    .Y(_12751_));
 sky130_fd_sc_hd__and2_2 _23031_ (.A(_12459_),
    .B(_12462_),
    .X(_12752_));
 sky130_fd_sc_hd__xnor2_2 _23032_ (.A(_12751_),
    .B(_12752_),
    .Y(_12753_));
 sky130_fd_sc_hd__nor2_2 _23033_ (.A(_11827_),
    .B(_12244_),
    .Y(_12755_));
 sky130_fd_sc_hd__and3_2 _23034_ (.A(_11783_),
    .B(_12242_),
    .C(_12755_),
    .X(_12756_));
 sky130_fd_sc_hd__a21oi_2 _23035_ (.A1(_11783_),
    .A2(_12242_),
    .B1(_12755_),
    .Y(_12757_));
 sky130_fd_sc_hd__nor2_2 _23036_ (.A(_12756_),
    .B(_12757_),
    .Y(_12758_));
 sky130_fd_sc_hd__buf_1 _23037_ (.A(_12477_),
    .X(_12759_));
 sky130_fd_sc_hd__nand2_2 _23038_ (.A(_11581_),
    .B(_12759_),
    .Y(_12760_));
 sky130_fd_sc_hd__xnor2_2 _23039_ (.A(_12758_),
    .B(_12760_),
    .Y(_12761_));
 sky130_fd_sc_hd__xnor2_2 _23040_ (.A(_12753_),
    .B(_12761_),
    .Y(_12762_));
 sky130_fd_sc_hd__and2b_2 _23041_ (.A_N(_12465_),
    .B(_12481_),
    .X(_12763_));
 sky130_fd_sc_hd__xnor2_2 _23042_ (.A(_12762_),
    .B(_12763_),
    .Y(_12764_));
 sky130_fd_sc_hd__and3_2 _23043_ (.A(_11374_),
    .B(_12471_),
    .C(_12759_),
    .X(_12766_));
 sky130_fd_sc_hd__nand2_2 _23044_ (.A(iY[6]),
    .B(iY[38]),
    .Y(_12767_));
 sky130_fd_sc_hd__or2_2 _23045_ (.A(iY[6]),
    .B(iY[38]),
    .X(_12768_));
 sky130_fd_sc_hd__nand2_2 _23046_ (.A(_12767_),
    .B(_12768_),
    .Y(_12769_));
 sky130_fd_sc_hd__or3_2 _23047_ (.A(_12236_),
    .B(_12237_),
    .C(_12474_),
    .X(_12770_));
 sky130_fd_sc_hd__o221ai_2 _23048_ (.A1(_12475_),
    .A2(_12474_),
    .B1(_12770_),
    .B2(_12239_),
    .C1(_12472_),
    .Y(_12771_));
 sky130_fd_sc_hd__xor2_2 _23049_ (.A(_12769_),
    .B(_12771_),
    .X(_12772_));
 sky130_fd_sc_hd__buf_1 _23050_ (.A(_12772_),
    .X(_12773_));
 sky130_fd_sc_hd__nor2_2 _23051_ (.A(_11577_),
    .B(_12773_),
    .Y(_12774_));
 sky130_fd_sc_hd__o21a_2 _23052_ (.A1(_12467_),
    .A2(_12766_),
    .B1(_12774_),
    .X(_12775_));
 sky130_fd_sc_hd__nor3_2 _23053_ (.A(_12467_),
    .B(_12766_),
    .C(_12774_),
    .Y(_12777_));
 sky130_fd_sc_hd__nor2_2 _23054_ (.A(_12775_),
    .B(_12777_),
    .Y(_12778_));
 sky130_fd_sc_hd__xor2_2 _23055_ (.A(_12764_),
    .B(_12778_),
    .X(_12779_));
 sky130_fd_sc_hd__and2b_2 _23056_ (.A_N(_12484_),
    .B(_12486_),
    .X(_12780_));
 sky130_fd_sc_hd__xnor2_2 _23057_ (.A(_12779_),
    .B(_12780_),
    .Y(_12781_));
 sky130_fd_sc_hd__or2_2 _23058_ (.A(_12488_),
    .B(_12781_),
    .X(_12782_));
 sky130_fd_sc_hd__nand2_2 _23059_ (.A(_12490_),
    .B(_12781_),
    .Y(_12783_));
 sky130_fd_sc_hd__nand2_2 _23060_ (.A(_12488_),
    .B(_12781_),
    .Y(_12784_));
 sky130_fd_sc_hd__o211a_2 _23061_ (.A1(_12490_),
    .A2(_12782_),
    .B1(_12783_),
    .C1(_12784_),
    .X(_12785_));
 sky130_fd_sc_hd__xnor2_2 _23062_ (.A(_12738_),
    .B(_12785_),
    .Y(_12786_));
 sky130_fd_sc_hd__xnor2_2 _23063_ (.A(_11923_),
    .B(_12786_),
    .Y(_12787_));
 sky130_fd_sc_hd__nand2_2 _23064_ (.A(_12522_),
    .B(_12525_),
    .Y(_12788_));
 sky130_fd_sc_hd__xor2_2 _23065_ (.A(_12787_),
    .B(_12788_),
    .X(_12789_));
 sky130_fd_sc_hd__a21oi_2 _23066_ (.A1(_12696_),
    .A2(_12697_),
    .B1(_12789_),
    .Y(_12790_));
 sky130_fd_sc_hd__and3_2 _23067_ (.A(_12696_),
    .B(_12697_),
    .C(_12789_),
    .X(_12791_));
 sky130_fd_sc_hd__nor2_2 _23068_ (.A(_12790_),
    .B(_12791_),
    .Y(_12792_));
 sky130_fd_sc_hd__nand2_2 _23069_ (.A(_12695_),
    .B(_12792_),
    .Y(_12793_));
 sky130_fd_sc_hd__or2_2 _23070_ (.A(_12695_),
    .B(_12792_),
    .X(_12794_));
 sky130_fd_sc_hd__nand2_2 _23071_ (.A(_12793_),
    .B(_12794_),
    .Y(_12795_));
 sky130_fd_sc_hd__a21o_2 _23072_ (.A1(_12292_),
    .A2(_12534_),
    .B1(_12536_),
    .X(_12796_));
 sky130_fd_sc_hd__xnor2_2 _23073_ (.A(_12795_),
    .B(_12796_),
    .Y(oO[38]));
 sky130_fd_sc_hd__inv_2 _23074_ (.A(_12286_),
    .Y(_12798_));
 sky130_fd_sc_hd__o211a_2 _23075_ (.A1(_12288_),
    .A2(_12289_),
    .B1(_12537_),
    .C1(_12798_),
    .X(_12799_));
 sky130_fd_sc_hd__or3b_2 _23076_ (.A(_12795_),
    .B(_12799_),
    .C_N(_12534_),
    .X(_12800_));
 sky130_fd_sc_hd__nand2_2 _23077_ (.A(_12783_),
    .B(_12784_),
    .Y(_12801_));
 sky130_fd_sc_hd__and2b_2 _23078_ (.A_N(_12780_),
    .B(_12779_),
    .X(_12802_));
 sky130_fd_sc_hd__or2b_2 _23079_ (.A(_12763_),
    .B_N(_12762_),
    .X(_12803_));
 sky130_fd_sc_hd__nand2_2 _23080_ (.A(_12764_),
    .B(_12778_),
    .Y(_12804_));
 sky130_fd_sc_hd__xor2_2 _23081_ (.A(iX[7]),
    .B(iX[39]),
    .X(_12805_));
 sky130_fd_sc_hd__a31oi_2 _23082_ (.A1(_12453_),
    .A2(_12742_),
    .A3(_12745_),
    .B1(_12740_),
    .Y(_12806_));
 sky130_fd_sc_hd__xor2_2 _23083_ (.A(_12805_),
    .B(_12806_),
    .X(_12808_));
 sky130_fd_sc_hd__nor3_2 _23084_ (.A(_11575_),
    .B(_12748_),
    .C(_12808_),
    .Y(_12809_));
 sky130_fd_sc_hd__nor2_2 _23085_ (.A(_12746_),
    .B(_12747_),
    .Y(_12810_));
 sky130_fd_sc_hd__xnor2_2 _23086_ (.A(_12805_),
    .B(_12806_),
    .Y(_12811_));
 sky130_fd_sc_hd__a22o_2 _23087_ (.A1(_11582_),
    .A2(_12810_),
    .B1(_12811_),
    .B2(_11379_),
    .X(_12812_));
 sky130_fd_sc_hd__or4b_2 _23088_ (.A(_11791_),
    .B(_12457_),
    .C(_12809_),
    .D_N(_12812_),
    .X(_12813_));
 sky130_fd_sc_hd__or3_2 _23089_ (.A(_11575_),
    .B(_12748_),
    .C(_12808_),
    .X(_12814_));
 sky130_fd_sc_hd__a22o_2 _23090_ (.A1(_12451_),
    .A2(_12460_),
    .B1(_12814_),
    .B2(_12812_),
    .X(_12815_));
 sky130_fd_sc_hd__buf_1 _23091_ (.A(_12810_),
    .X(_12816_));
 sky130_fd_sc_hd__and3_2 _23092_ (.A(_11380_),
    .B(_12739_),
    .C(_12816_),
    .X(_12817_));
 sky130_fd_sc_hd__a21o_2 _23093_ (.A1(_12749_),
    .A2(_12750_),
    .B1(_12817_),
    .X(_12819_));
 sky130_fd_sc_hd__nand3_2 _23094_ (.A(_12813_),
    .B(_12815_),
    .C(_12819_),
    .Y(_12820_));
 sky130_fd_sc_hd__a21o_2 _23095_ (.A1(_12813_),
    .A2(_12815_),
    .B1(_12819_),
    .X(_12821_));
 sky130_fd_sc_hd__nand2_2 _23096_ (.A(_11829_),
    .B(_11842_),
    .Y(_12822_));
 sky130_fd_sc_hd__nand2_2 _23097_ (.A(_12225_),
    .B(_12241_),
    .Y(_12823_));
 sky130_fd_sc_hd__nor2_2 _23098_ (.A(_12822_),
    .B(_12823_),
    .Y(_12824_));
 sky130_fd_sc_hd__o22a_2 _23099_ (.A1(_12244_),
    .A2(_12223_),
    .B1(_12248_),
    .B2(_11827_),
    .X(_12825_));
 sky130_fd_sc_hd__nor2_2 _23100_ (.A(_12824_),
    .B(_12825_),
    .Y(_12826_));
 sky130_fd_sc_hd__buf_1 _23101_ (.A(_11783_),
    .X(_12827_));
 sky130_fd_sc_hd__nand2_2 _23102_ (.A(_12827_),
    .B(_12477_),
    .Y(_12828_));
 sky130_fd_sc_hd__xnor2_2 _23103_ (.A(_12826_),
    .B(_12828_),
    .Y(_12830_));
 sky130_fd_sc_hd__nand3_2 _23104_ (.A(_12820_),
    .B(_12821_),
    .C(_12830_),
    .Y(_12831_));
 sky130_fd_sc_hd__a21o_2 _23105_ (.A1(_12820_),
    .A2(_12821_),
    .B1(_12830_),
    .X(_12832_));
 sky130_fd_sc_hd__nand2_2 _23106_ (.A(_12751_),
    .B(_12752_),
    .Y(_12833_));
 sky130_fd_sc_hd__nor2_2 _23107_ (.A(_12751_),
    .B(_12752_),
    .Y(_12834_));
 sky130_fd_sc_hd__a21o_2 _23108_ (.A1(_12833_),
    .A2(_12761_),
    .B1(_12834_),
    .X(_12835_));
 sky130_fd_sc_hd__and3_2 _23109_ (.A(_12831_),
    .B(_12832_),
    .C(_12835_),
    .X(_12836_));
 sky130_fd_sc_hd__a21oi_2 _23110_ (.A1(_12831_),
    .A2(_12832_),
    .B1(_12835_),
    .Y(_12837_));
 sky130_fd_sc_hd__buf_1 _23111_ (.A(_11581_),
    .X(_12838_));
 sky130_fd_sc_hd__a31o_2 _23112_ (.A1(_12838_),
    .A2(_12759_),
    .A3(_12758_),
    .B1(_12756_),
    .X(_12839_));
 sky130_fd_sc_hd__nand2_2 _23113_ (.A(iY[7]),
    .B(iY[39]),
    .Y(_12841_));
 sky130_fd_sc_hd__or2_2 _23114_ (.A(iY[7]),
    .B(iY[39]),
    .X(_12842_));
 sky130_fd_sc_hd__nand2_2 _23115_ (.A(_12841_),
    .B(_12842_),
    .Y(_12843_));
 sky130_fd_sc_hd__a21boi_2 _23116_ (.A1(_12768_),
    .A2(_12771_),
    .B1_N(_12767_),
    .Y(_12844_));
 sky130_fd_sc_hd__xor2_2 _23117_ (.A(_12843_),
    .B(_12844_),
    .X(_12845_));
 sky130_fd_sc_hd__buf_1 _23118_ (.A(_12845_),
    .X(_12846_));
 sky130_fd_sc_hd__and3_2 _23119_ (.A(_11581_),
    .B(_12774_),
    .C(_12846_),
    .X(_12847_));
 sky130_fd_sc_hd__buf_1 _23120_ (.A(_12773_),
    .X(_12848_));
 sky130_fd_sc_hd__xnor2_2 _23121_ (.A(_12843_),
    .B(_12844_),
    .Y(_12849_));
 sky130_fd_sc_hd__buf_1 _23122_ (.A(_12849_),
    .X(_12850_));
 sky130_fd_sc_hd__buf_1 _23123_ (.A(_12850_),
    .X(_12852_));
 sky130_fd_sc_hd__o22a_2 _23124_ (.A1(_11570_),
    .A2(_12848_),
    .B1(_12852_),
    .B2(_11577_),
    .X(_12853_));
 sky130_fd_sc_hd__or2_2 _23125_ (.A(_12847_),
    .B(_12853_),
    .X(_12854_));
 sky130_fd_sc_hd__xor2_2 _23126_ (.A(_12839_),
    .B(_12854_),
    .X(_12855_));
 sky130_fd_sc_hd__nor3_2 _23127_ (.A(_12836_),
    .B(_12837_),
    .C(_12855_),
    .Y(_12856_));
 sky130_fd_sc_hd__o21a_2 _23128_ (.A1(_12836_),
    .A2(_12837_),
    .B1(_12855_),
    .X(_12857_));
 sky130_fd_sc_hd__a211o_2 _23129_ (.A1(_12803_),
    .A2(_12804_),
    .B1(_12856_),
    .C1(_12857_),
    .X(_12858_));
 sky130_fd_sc_hd__o211ai_2 _23130_ (.A1(_12856_),
    .A2(_12857_),
    .B1(_12803_),
    .C1(_12804_),
    .Y(_12859_));
 sky130_fd_sc_hd__nand3_2 _23131_ (.A(_12775_),
    .B(_12858_),
    .C(_12859_),
    .Y(_12860_));
 sky130_fd_sc_hd__a21o_2 _23132_ (.A1(_12858_),
    .A2(_12859_),
    .B1(_12775_),
    .X(_12861_));
 sky130_fd_sc_hd__and3_2 _23133_ (.A(_12802_),
    .B(_12860_),
    .C(_12861_),
    .X(_12863_));
 sky130_fd_sc_hd__a21oi_2 _23134_ (.A1(_12860_),
    .A2(_12861_),
    .B1(_12802_),
    .Y(_12864_));
 sky130_fd_sc_hd__or3_2 _23135_ (.A(_12801_),
    .B(_12863_),
    .C(_12864_),
    .X(_12865_));
 sky130_fd_sc_hd__o21ai_2 _23136_ (.A1(_12863_),
    .A2(_12864_),
    .B1(_12801_),
    .Y(_12866_));
 sky130_fd_sc_hd__and3b_2 _23137_ (.A_N(_12717_),
    .B(_12719_),
    .C(_12724_),
    .X(_12867_));
 sky130_fd_sc_hd__and4_2 _23138_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[36]),
    .D(iX[37]),
    .X(_12868_));
 sky130_fd_sc_hd__a22oi_2 _23139_ (.A1(iY[35]),
    .A2(iX[36]),
    .B1(iX[37]),
    .B2(iY[34]),
    .Y(_12869_));
 sky130_fd_sc_hd__nand2_2 _23140_ (.A(iY[33]),
    .B(iX[38]),
    .Y(_12870_));
 sky130_fd_sc_hd__or3_2 _23141_ (.A(_12868_),
    .B(_12869_),
    .C(_12870_),
    .X(_12871_));
 sky130_fd_sc_hd__o21ai_2 _23142_ (.A1(_12868_),
    .A2(_12869_),
    .B1(_12870_),
    .Y(_12872_));
 sky130_fd_sc_hd__o21bai_2 _23143_ (.A1(_12701_),
    .A2(_12702_),
    .B1_N(_12700_),
    .Y(_12874_));
 sky130_fd_sc_hd__nand3_2 _23144_ (.A(_12871_),
    .B(_12872_),
    .C(_12874_),
    .Y(_12875_));
 sky130_fd_sc_hd__a21o_2 _23145_ (.A1(_12871_),
    .A2(_12872_),
    .B1(_12874_),
    .X(_12876_));
 sky130_fd_sc_hd__and4_2 _23146_ (.A(iY[32]),
    .B(iX[35]),
    .C(iY[36]),
    .D(iX[39]),
    .X(_12877_));
 sky130_fd_sc_hd__a22o_2 _23147_ (.A1(iX[35]),
    .A2(iY[36]),
    .B1(iX[39]),
    .B2(iY[32]),
    .X(_12878_));
 sky130_fd_sc_hd__and2b_2 _23148_ (.A_N(_12877_),
    .B(_12878_),
    .X(_12879_));
 sky130_fd_sc_hd__nand2_2 _23149_ (.A(iX[34]),
    .B(iY[37]),
    .Y(_12880_));
 sky130_fd_sc_hd__xnor2_2 _23150_ (.A(_12879_),
    .B(_12880_),
    .Y(_12881_));
 sky130_fd_sc_hd__nand3_2 _23151_ (.A(_12875_),
    .B(_12876_),
    .C(_12881_),
    .Y(_12882_));
 sky130_fd_sc_hd__a21o_2 _23152_ (.A1(_12875_),
    .A2(_12876_),
    .B1(_12881_),
    .X(_12883_));
 sky130_fd_sc_hd__a21bo_2 _23153_ (.A1(_12707_),
    .A2(_12713_),
    .B1_N(_12706_),
    .X(_12885_));
 sky130_fd_sc_hd__nand3_2 _23154_ (.A(_12882_),
    .B(_12883_),
    .C(_12885_),
    .Y(_12886_));
 sky130_fd_sc_hd__a21o_2 _23155_ (.A1(_12882_),
    .A2(_12883_),
    .B1(_12885_),
    .X(_12887_));
 sky130_fd_sc_hd__and4_2 _23156_ (.A(iX[33]),
    .B(iX[32]),
    .C(iY[38]),
    .D(iY[39]),
    .X(_12888_));
 sky130_fd_sc_hd__a22oi_2 _23157_ (.A1(iX[33]),
    .A2(iY[38]),
    .B1(iY[39]),
    .B2(iX[32]),
    .Y(_12889_));
 sky130_fd_sc_hd__or2_2 _23158_ (.A(_12888_),
    .B(_12889_),
    .X(_12890_));
 sky130_fd_sc_hd__a32o_2 _23159_ (.A1(iX[33]),
    .A2(iY[37]),
    .A3(_12709_),
    .B1(_12708_),
    .B2(iY[36]),
    .X(_12891_));
 sky130_fd_sc_hd__and2b_2 _23160_ (.A_N(_12890_),
    .B(_12891_),
    .X(_12892_));
 sky130_fd_sc_hd__and2b_2 _23161_ (.A_N(_12891_),
    .B(_12890_),
    .X(_12893_));
 sky130_fd_sc_hd__nor2_2 _23162_ (.A(_12892_),
    .B(_12893_),
    .Y(_12894_));
 sky130_fd_sc_hd__nand3_2 _23163_ (.A(_12886_),
    .B(_12887_),
    .C(_12894_),
    .Y(_12896_));
 sky130_fd_sc_hd__a21o_2 _23164_ (.A1(_12886_),
    .A2(_12887_),
    .B1(_12894_),
    .X(_12897_));
 sky130_fd_sc_hd__o211ai_2 _23165_ (.A1(_12717_),
    .A2(_12867_),
    .B1(_12896_),
    .C1(_12897_),
    .Y(_12898_));
 sky130_fd_sc_hd__a211o_2 _23166_ (.A1(_12896_),
    .A2(_12897_),
    .B1(_12717_),
    .C1(_12867_),
    .X(_12899_));
 sky130_fd_sc_hd__nand3_2 _23167_ (.A(_12722_),
    .B(_12898_),
    .C(_12899_),
    .Y(_12900_));
 sky130_fd_sc_hd__a21o_2 _23168_ (.A1(_12898_),
    .A2(_12899_),
    .B1(_12722_),
    .X(_12901_));
 sky130_fd_sc_hd__nand3b_2 _23169_ (.A_N(_12727_),
    .B(_12900_),
    .C(_12901_),
    .Y(_12902_));
 sky130_fd_sc_hd__a21bo_2 _23170_ (.A1(_12900_),
    .A2(_12901_),
    .B1_N(_12727_),
    .X(_12903_));
 sky130_fd_sc_hd__nand2_2 _23171_ (.A(_12902_),
    .B(_12903_),
    .Y(_12904_));
 sky130_fd_sc_hd__inv_2 _23172_ (.A(_12729_),
    .Y(_12905_));
 sky130_fd_sc_hd__and2_2 _23173_ (.A(_12905_),
    .B(_12733_),
    .X(_12907_));
 sky130_fd_sc_hd__xnor2_2 _23174_ (.A(_12904_),
    .B(_12907_),
    .Y(_12908_));
 sky130_fd_sc_hd__and2b_2 _23175_ (.A_N(_12908_),
    .B(_12736_),
    .X(_12909_));
 sky130_fd_sc_hd__and2b_2 _23176_ (.A_N(_12736_),
    .B(_12908_),
    .X(_12910_));
 sky130_fd_sc_hd__nor2_2 _23177_ (.A(_12909_),
    .B(_12910_),
    .Y(_12911_));
 sky130_fd_sc_hd__a21o_2 _23178_ (.A1(_12865_),
    .A2(_12866_),
    .B1(_12911_),
    .X(_12912_));
 sky130_fd_sc_hd__nand3_2 _23179_ (.A(_12911_),
    .B(_12865_),
    .C(_12866_),
    .Y(_12913_));
 sky130_fd_sc_hd__nand2_2 _23180_ (.A(_12912_),
    .B(_12913_),
    .Y(_12914_));
 sky130_fd_sc_hd__xnor2_2 _23181_ (.A(_12327_),
    .B(_12914_),
    .Y(_12915_));
 sky130_fd_sc_hd__and2b_2 _23182_ (.A_N(_12738_),
    .B(_12785_),
    .X(_12916_));
 sky130_fd_sc_hd__a21o_2 _23183_ (.A1(_11923_),
    .A2(_12786_),
    .B1(_12916_),
    .X(_12918_));
 sky130_fd_sc_hd__xnor2_2 _23184_ (.A(_12915_),
    .B(_12918_),
    .Y(_12919_));
 sky130_fd_sc_hd__and2b_2 _23185_ (.A_N(_12787_),
    .B(_12788_),
    .X(_12920_));
 sky130_fd_sc_hd__nor2_2 _23186_ (.A(_12920_),
    .B(_12790_),
    .Y(_12921_));
 sky130_fd_sc_hd__xnor2_2 _23187_ (.A(_12919_),
    .B(_12921_),
    .Y(_12922_));
 sky130_fd_sc_hd__and2b_2 _23188_ (.A_N(_12682_),
    .B(_12683_),
    .X(_12923_));
 sky130_fd_sc_hd__and2b_2 _23189_ (.A_N(_12607_),
    .B(_12606_),
    .X(_12924_));
 sky130_fd_sc_hd__a21oi_2 _23190_ (.A1(_12599_),
    .A2(_12608_),
    .B1(_12924_),
    .Y(_12925_));
 sky130_fd_sc_hd__and4_2 _23191_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[26]),
    .D(iX[27]),
    .X(_12926_));
 sky130_fd_sc_hd__a22oi_2 _23192_ (.A1(iY[13]),
    .A2(iX[26]),
    .B1(iX[27]),
    .B2(iY[12]),
    .Y(_12927_));
 sky130_fd_sc_hd__nor2_2 _23193_ (.A(_12926_),
    .B(_12927_),
    .Y(_12929_));
 sky130_fd_sc_hd__nand2_2 _23194_ (.A(iY[14]),
    .B(iX[25]),
    .Y(_12930_));
 sky130_fd_sc_hd__xnor2_2 _23195_ (.A(_12929_),
    .B(_12930_),
    .Y(_12931_));
 sky130_fd_sc_hd__and2_2 _23196_ (.A(iY[10]),
    .B(iX[30]),
    .X(_12932_));
 sky130_fd_sc_hd__a22oi_2 _23197_ (.A1(iY[10]),
    .A2(iX[29]),
    .B1(iX[30]),
    .B2(iY[9]),
    .Y(_12933_));
 sky130_fd_sc_hd__a21o_2 _23198_ (.A1(_12602_),
    .A2(_12932_),
    .B1(_12933_),
    .X(_12934_));
 sky130_fd_sc_hd__nand2_2 _23199_ (.A(iY[11]),
    .B(iX[28]),
    .Y(_12935_));
 sky130_fd_sc_hd__xor2_2 _23200_ (.A(_12934_),
    .B(_12935_),
    .X(_12936_));
 sky130_fd_sc_hd__o21ba_2 _23201_ (.A1(_12603_),
    .A2(_12605_),
    .B1_N(_12601_),
    .X(_12937_));
 sky130_fd_sc_hd__xnor2_2 _23202_ (.A(_12936_),
    .B(_12937_),
    .Y(_12938_));
 sky130_fd_sc_hd__xnor2_2 _23203_ (.A(_12931_),
    .B(_12938_),
    .Y(_12940_));
 sky130_fd_sc_hd__or2_2 _23204_ (.A(_12591_),
    .B(_12940_),
    .X(_12941_));
 sky130_fd_sc_hd__nand2_2 _23205_ (.A(_12591_),
    .B(_12940_),
    .Y(_12942_));
 sky130_fd_sc_hd__and2_2 _23206_ (.A(_12941_),
    .B(_12942_),
    .X(_12943_));
 sky130_fd_sc_hd__xnor2_2 _23207_ (.A(_12925_),
    .B(_12943_),
    .Y(_12944_));
 sky130_fd_sc_hd__and3b_2 _23208_ (.A_N(_12586_),
    .B(_12944_),
    .C(_12050_),
    .X(_12945_));
 sky130_fd_sc_hd__o21ba_2 _23209_ (.A1(_12296_),
    .A2(_12586_),
    .B1_N(_12944_),
    .X(_12946_));
 sky130_fd_sc_hd__or2_2 _23210_ (.A(_12945_),
    .B(_12946_),
    .X(_12947_));
 sky130_fd_sc_hd__xnor2_2 _23211_ (.A(_12616_),
    .B(_12947_),
    .Y(_12948_));
 sky130_fd_sc_hd__inv_2 _23212_ (.A(_12576_),
    .Y(_12949_));
 sky130_fd_sc_hd__and4_2 _23213_ (.A(iX[17]),
    .B(iX[18]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_12951_));
 sky130_fd_sc_hd__a22oi_2 _23214_ (.A1(iX[18]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[17]),
    .Y(_12952_));
 sky130_fd_sc_hd__nor2_2 _23215_ (.A(_12951_),
    .B(_12952_),
    .Y(_12953_));
 sky130_fd_sc_hd__nand2_2 _23216_ (.A(iX[16]),
    .B(iY[23]),
    .Y(_12954_));
 sky130_fd_sc_hd__xnor2_2 _23217_ (.A(_12953_),
    .B(_12954_),
    .Y(_12955_));
 sky130_fd_sc_hd__and4_2 _23218_ (.A(iY[18]),
    .B(iY[19]),
    .C(iX[20]),
    .D(iX[21]),
    .X(_12956_));
 sky130_fd_sc_hd__a22oi_2 _23219_ (.A1(iY[19]),
    .A2(iX[20]),
    .B1(iX[21]),
    .B2(iY[18]),
    .Y(_12957_));
 sky130_fd_sc_hd__nor2_2 _23220_ (.A(_12956_),
    .B(_12957_),
    .Y(_12958_));
 sky130_fd_sc_hd__nand2_2 _23221_ (.A(iX[19]),
    .B(iY[20]),
    .Y(_12959_));
 sky130_fd_sc_hd__xnor2_2 _23222_ (.A(_12958_),
    .B(_12959_),
    .Y(_12960_));
 sky130_fd_sc_hd__o21ba_2 _23223_ (.A1(_12552_),
    .A2(_12554_),
    .B1_N(_12551_),
    .X(_12962_));
 sky130_fd_sc_hd__xnor2_2 _23224_ (.A(_12960_),
    .B(_12962_),
    .Y(_12963_));
 sky130_fd_sc_hd__and2_2 _23225_ (.A(_12955_),
    .B(_12963_),
    .X(_12964_));
 sky130_fd_sc_hd__nor2_2 _23226_ (.A(_12955_),
    .B(_12963_),
    .Y(_12965_));
 sky130_fd_sc_hd__or2_2 _23227_ (.A(_12964_),
    .B(_12965_),
    .X(_12966_));
 sky130_fd_sc_hd__or3_2 _23228_ (.A(_12564_),
    .B(_12569_),
    .C(_12570_),
    .X(_12967_));
 sky130_fd_sc_hd__o21ba_2 _23229_ (.A1(_12596_),
    .A2(_12598_),
    .B1_N(_12595_),
    .X(_12968_));
 sky130_fd_sc_hd__and4_2 _23230_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[23]),
    .D(iX[24]),
    .X(_12969_));
 sky130_fd_sc_hd__a22oi_2 _23231_ (.A1(iY[16]),
    .A2(iX[23]),
    .B1(iX[24]),
    .B2(iY[15]),
    .Y(_12970_));
 sky130_fd_sc_hd__nand2_2 _23232_ (.A(iY[17]),
    .B(iX[22]),
    .Y(_12971_));
 sky130_fd_sc_hd__o21a_2 _23233_ (.A1(_12969_),
    .A2(_12970_),
    .B1(_12971_),
    .X(_12973_));
 sky130_fd_sc_hd__nor3_2 _23234_ (.A(_12969_),
    .B(_12970_),
    .C(_12971_),
    .Y(_12974_));
 sky130_fd_sc_hd__nor2_2 _23235_ (.A(_12973_),
    .B(_12974_),
    .Y(_12975_));
 sky130_fd_sc_hd__xnor2_2 _23236_ (.A(_12968_),
    .B(_12975_),
    .Y(_12976_));
 sky130_fd_sc_hd__o21ai_2 _23237_ (.A1(_12565_),
    .A2(_12570_),
    .B1(_12976_),
    .Y(_12977_));
 sky130_fd_sc_hd__or3_2 _23238_ (.A(_12565_),
    .B(_12570_),
    .C(_12976_),
    .X(_12978_));
 sky130_fd_sc_hd__nand2_2 _23239_ (.A(_12977_),
    .B(_12978_),
    .Y(_12979_));
 sky130_fd_sc_hd__a21oi_2 _23240_ (.A1(_12967_),
    .A2(_12573_),
    .B1(_12979_),
    .Y(_12980_));
 sky130_fd_sc_hd__and3_2 _23241_ (.A(_12967_),
    .B(_12573_),
    .C(_12979_),
    .X(_12981_));
 sky130_fd_sc_hd__or3_2 _23242_ (.A(_12966_),
    .B(_12980_),
    .C(_12981_),
    .X(_12982_));
 sky130_fd_sc_hd__o21ai_2 _23243_ (.A1(_12980_),
    .A2(_12981_),
    .B1(_12966_),
    .Y(_12984_));
 sky130_fd_sc_hd__nand2_2 _23244_ (.A(_12982_),
    .B(_12984_),
    .Y(_12985_));
 sky130_fd_sc_hd__a21oi_2 _23245_ (.A1(_12610_),
    .A2(_12614_),
    .B1(_12985_),
    .Y(_12986_));
 sky130_fd_sc_hd__and3_2 _23246_ (.A(_12610_),
    .B(_12614_),
    .C(_12985_),
    .X(_12987_));
 sky130_fd_sc_hd__a211o_2 _23247_ (.A1(_12949_),
    .A2(_12579_),
    .B1(_12986_),
    .C1(_12987_),
    .X(_12988_));
 sky130_fd_sc_hd__o211ai_2 _23248_ (.A1(_12986_),
    .A2(_12987_),
    .B1(_12949_),
    .C1(_12579_),
    .Y(_12989_));
 sky130_fd_sc_hd__nand3_2 _23249_ (.A(_12948_),
    .B(_12988_),
    .C(_12989_),
    .Y(_12990_));
 sky130_fd_sc_hd__a21o_2 _23250_ (.A1(_12988_),
    .A2(_12989_),
    .B1(_12948_),
    .X(_12991_));
 sky130_fd_sc_hd__nand2_2 _23251_ (.A(_12990_),
    .B(_12991_),
    .Y(_12992_));
 sky130_fd_sc_hd__a21oi_2 _23252_ (.A1(_12618_),
    .A2(_12623_),
    .B1(_12992_),
    .Y(_12993_));
 sky130_fd_sc_hd__and3_2 _23253_ (.A(_12618_),
    .B(_12623_),
    .C(_12992_),
    .X(_12995_));
 sky130_fd_sc_hd__inv_2 _23254_ (.A(_12668_),
    .Y(_12996_));
 sky130_fd_sc_hd__or2b_2 _23255_ (.A(_12634_),
    .B_N(_12632_),
    .X(_12997_));
 sky130_fd_sc_hd__and4_2 _23256_ (.A(iX[11]),
    .B(iX[12]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_12998_));
 sky130_fd_sc_hd__a22oi_2 _23257_ (.A1(iX[12]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[11]),
    .Y(_12999_));
 sky130_fd_sc_hd__nor2_2 _23258_ (.A(_12998_),
    .B(_12999_),
    .Y(_13000_));
 sky130_fd_sc_hd__nand2_2 _23259_ (.A(iX[10]),
    .B(iY[29]),
    .Y(_13001_));
 sky130_fd_sc_hd__xnor2_2 _23260_ (.A(_13000_),
    .B(_13001_),
    .Y(_13002_));
 sky130_fd_sc_hd__o21ba_2 _23261_ (.A1(_12629_),
    .A2(_12631_),
    .B1_N(_12628_),
    .X(_13003_));
 sky130_fd_sc_hd__xnor2_2 _23262_ (.A(_13002_),
    .B(_13003_),
    .Y(_13004_));
 sky130_fd_sc_hd__and2_2 _23263_ (.A(iX[9]),
    .B(iY[30]),
    .X(_13006_));
 sky130_fd_sc_hd__or2_2 _23264_ (.A(_13004_),
    .B(_13006_),
    .X(_13007_));
 sky130_fd_sc_hd__nand2_2 _23265_ (.A(_13004_),
    .B(_13006_),
    .Y(_13008_));
 sky130_fd_sc_hd__nand2_2 _23266_ (.A(_13007_),
    .B(_13008_),
    .Y(_13009_));
 sky130_fd_sc_hd__a21oi_2 _23267_ (.A1(_12997_),
    .A2(_12638_),
    .B1(_13009_),
    .Y(_13010_));
 sky130_fd_sc_hd__and3_2 _23268_ (.A(_12997_),
    .B(_12638_),
    .C(_13009_),
    .X(_13011_));
 sky130_fd_sc_hd__nor2_2 _23269_ (.A(_13010_),
    .B(_13011_),
    .Y(_13012_));
 sky130_fd_sc_hd__nand2_2 _23270_ (.A(iX[8]),
    .B(iY[31]),
    .Y(_13013_));
 sky130_fd_sc_hd__xnor2_2 _23271_ (.A(_13012_),
    .B(_13013_),
    .Y(_13014_));
 sky130_fd_sc_hd__or2b_2 _23272_ (.A(_12653_),
    .B_N(_12659_),
    .X(_13015_));
 sky130_fd_sc_hd__or2b_2 _23273_ (.A(_12652_),
    .B_N(_12660_),
    .X(_13017_));
 sky130_fd_sc_hd__and2b_2 _23274_ (.A_N(_12557_),
    .B(_12555_),
    .X(_13018_));
 sky130_fd_sc_hd__o21ba_2 _23275_ (.A1(_12656_),
    .A2(_12658_),
    .B1_N(_12654_),
    .X(_13019_));
 sky130_fd_sc_hd__o21ba_2 _23276_ (.A1(_12547_),
    .A2(_12549_),
    .B1_N(_12546_),
    .X(_13020_));
 sky130_fd_sc_hd__and4_2 _23277_ (.A(iX[14]),
    .B(iX[15]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_13021_));
 sky130_fd_sc_hd__a22oi_2 _23278_ (.A1(iX[15]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[14]),
    .Y(_13022_));
 sky130_fd_sc_hd__nor2_2 _23279_ (.A(_13021_),
    .B(_13022_),
    .Y(_13023_));
 sky130_fd_sc_hd__nand2_2 _23280_ (.A(iX[13]),
    .B(iY[26]),
    .Y(_13024_));
 sky130_fd_sc_hd__xnor2_2 _23281_ (.A(_13023_),
    .B(_13024_),
    .Y(_13025_));
 sky130_fd_sc_hd__xnor2_2 _23282_ (.A(_13020_),
    .B(_13025_),
    .Y(_13026_));
 sky130_fd_sc_hd__xnor2_2 _23283_ (.A(_13019_),
    .B(_13026_),
    .Y(_13028_));
 sky130_fd_sc_hd__o21a_2 _23284_ (.A1(_13018_),
    .A2(_12559_),
    .B1(_13028_),
    .X(_13029_));
 sky130_fd_sc_hd__nor3_2 _23285_ (.A(_13018_),
    .B(_12559_),
    .C(_13028_),
    .Y(_13030_));
 sky130_fd_sc_hd__a211oi_2 _23286_ (.A1(_13015_),
    .A2(_13017_),
    .B1(_13029_),
    .C1(_13030_),
    .Y(_13031_));
 sky130_fd_sc_hd__o211a_2 _23287_ (.A1(_13029_),
    .A2(_13030_),
    .B1(_13015_),
    .C1(_13017_),
    .X(_13032_));
 sky130_fd_sc_hd__nor2_2 _23288_ (.A(_12662_),
    .B(_12664_),
    .Y(_13033_));
 sky130_fd_sc_hd__or3_2 _23289_ (.A(_13031_),
    .B(_13032_),
    .C(_13033_),
    .X(_13034_));
 sky130_fd_sc_hd__o21ai_2 _23290_ (.A1(_13031_),
    .A2(_13032_),
    .B1(_13033_),
    .Y(_13035_));
 sky130_fd_sc_hd__and3_2 _23291_ (.A(_13014_),
    .B(_13034_),
    .C(_13035_),
    .X(_13036_));
 sky130_fd_sc_hd__a21oi_2 _23292_ (.A1(_13034_),
    .A2(_13035_),
    .B1(_13014_),
    .Y(_13037_));
 sky130_fd_sc_hd__nor2_2 _23293_ (.A(_13036_),
    .B(_13037_),
    .Y(_13039_));
 sky130_fd_sc_hd__o21ai_2 _23294_ (.A1(_12582_),
    .A2(_12584_),
    .B1(_13039_),
    .Y(_13040_));
 sky130_fd_sc_hd__or3_2 _23295_ (.A(_12582_),
    .B(_12584_),
    .C(_13039_),
    .X(_13041_));
 sky130_fd_sc_hd__o211ai_2 _23296_ (.A1(_12996_),
    .A2(_12670_),
    .B1(_13040_),
    .C1(_13041_),
    .Y(_13042_));
 sky130_fd_sc_hd__a211o_2 _23297_ (.A1(_13040_),
    .A2(_13041_),
    .B1(_12996_),
    .C1(_12670_),
    .X(_13043_));
 sky130_fd_sc_hd__or4bb_2 _23298_ (.A(_12993_),
    .B(_12995_),
    .C_N(_13042_),
    .D_N(_13043_),
    .X(_13044_));
 sky130_fd_sc_hd__a2bb2o_2 _23299_ (.A1_N(_12993_),
    .A2_N(_12995_),
    .B1(_13042_),
    .B2(_13043_),
    .X(_13045_));
 sky130_fd_sc_hd__nand2_2 _23300_ (.A(_12625_),
    .B(_12678_),
    .Y(_13046_));
 sky130_fd_sc_hd__and3_2 _23301_ (.A(_13044_),
    .B(_13045_),
    .C(_13046_),
    .X(_13047_));
 sky130_fd_sc_hd__a21oi_2 _23302_ (.A1(_13044_),
    .A2(_13045_),
    .B1(_13046_),
    .Y(_13048_));
 sky130_fd_sc_hd__a211oi_2 _23303_ (.A1(_12673_),
    .A2(_12675_),
    .B1(_13047_),
    .C1(_13048_),
    .Y(_13050_));
 sky130_fd_sc_hd__o211a_2 _23304_ (.A1(_13047_),
    .A2(_13048_),
    .B1(_12673_),
    .C1(_12675_),
    .X(_13051_));
 sky130_fd_sc_hd__nor2_2 _23305_ (.A(_13050_),
    .B(_13051_),
    .Y(_13052_));
 sky130_fd_sc_hd__o21a_2 _23306_ (.A1(_12680_),
    .A2(_12923_),
    .B1(_13052_),
    .X(_13053_));
 sky130_fd_sc_hd__nor3_2 _23307_ (.A(_12680_),
    .B(_12923_),
    .C(_13052_),
    .Y(_13054_));
 sky130_fd_sc_hd__a211oi_2 _23308_ (.A1(_12641_),
    .A2(_12647_),
    .B1(_13053_),
    .C1(_13054_),
    .Y(_13055_));
 sky130_fd_sc_hd__o211a_2 _23309_ (.A1(_13053_),
    .A2(_13054_),
    .B1(_12641_),
    .C1(_12647_),
    .X(_13056_));
 sky130_fd_sc_hd__or2b_2 _23310_ (.A(_12687_),
    .B_N(_12689_),
    .X(_13057_));
 sky130_fd_sc_hd__o211a_2 _23311_ (.A1(_13055_),
    .A2(_13056_),
    .B1(_12685_),
    .C1(_13057_),
    .X(_13058_));
 sky130_fd_sc_hd__a211oi_2 _23312_ (.A1(_12685_),
    .A2(_13057_),
    .B1(_13055_),
    .C1(_13056_),
    .Y(_13059_));
 sky130_fd_sc_hd__or2_2 _23313_ (.A(_13058_),
    .B(_13059_),
    .X(_13061_));
 sky130_fd_sc_hd__inv_2 _23314_ (.A(_12693_),
    .Y(_13062_));
 sky130_fd_sc_hd__a21oi_2 _23315_ (.A1(_13062_),
    .A2(_12694_),
    .B1(_12691_),
    .Y(_13063_));
 sky130_fd_sc_hd__xnor2_2 _23316_ (.A(_13061_),
    .B(_13063_),
    .Y(_13064_));
 sky130_fd_sc_hd__nor2_2 _23317_ (.A(_12922_),
    .B(_13064_),
    .Y(_13065_));
 sky130_fd_sc_hd__and2_2 _23318_ (.A(_12922_),
    .B(_13064_),
    .X(_13066_));
 sky130_fd_sc_hd__or2_2 _23319_ (.A(_13065_),
    .B(_13066_),
    .X(_13067_));
 sky130_fd_sc_hd__a21oi_2 _23320_ (.A1(_12793_),
    .A2(_12800_),
    .B1(_13067_),
    .Y(_13068_));
 sky130_fd_sc_hd__and3_2 _23321_ (.A(_12793_),
    .B(_12800_),
    .C(_13067_),
    .X(_13069_));
 sky130_fd_sc_hd__nor2_2 _23322_ (.A(_13068_),
    .B(_13069_),
    .Y(oO[39]));
 sky130_fd_sc_hd__inv_2 _23323_ (.A(_13065_),
    .Y(_13071_));
 sky130_fd_sc_hd__a21o_2 _23324_ (.A1(_12793_),
    .A2(_12800_),
    .B1(_13067_),
    .X(_13072_));
 sky130_fd_sc_hd__nand2_2 _23325_ (.A(_13071_),
    .B(_13072_),
    .Y(_13073_));
 sky130_fd_sc_hd__inv_2 _23326_ (.A(_13044_),
    .Y(_13074_));
 sky130_fd_sc_hd__or3b_2 _23327_ (.A(_12945_),
    .B(_12946_),
    .C_N(_12616_),
    .X(_13075_));
 sky130_fd_sc_hd__inv_2 _23328_ (.A(_12945_),
    .Y(_13076_));
 sky130_fd_sc_hd__and4_2 _23329_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[27]),
    .D(iX[28]),
    .X(_13077_));
 sky130_fd_sc_hd__a22oi_2 _23330_ (.A1(iY[13]),
    .A2(iX[27]),
    .B1(iX[28]),
    .B2(iY[12]),
    .Y(_13078_));
 sky130_fd_sc_hd__or2_2 _23331_ (.A(_13077_),
    .B(_13078_),
    .X(_13079_));
 sky130_fd_sc_hd__nand2_2 _23332_ (.A(iY[14]),
    .B(iX[26]),
    .Y(_13080_));
 sky130_fd_sc_hd__nor2_2 _23333_ (.A(_13079_),
    .B(_13080_),
    .Y(_13082_));
 sky130_fd_sc_hd__and2_2 _23334_ (.A(_13079_),
    .B(_13080_),
    .X(_13083_));
 sky130_fd_sc_hd__nor2_2 _23335_ (.A(_13082_),
    .B(_13083_),
    .Y(_13084_));
 sky130_fd_sc_hd__inv_2 _23336_ (.A(_13084_),
    .Y(_13085_));
 sky130_fd_sc_hd__a21o_2 _23337_ (.A1(iY[9]),
    .A2(iX[31]),
    .B1(_12932_),
    .X(_13086_));
 sky130_fd_sc_hd__and3_2 _23338_ (.A(iY[9]),
    .B(iX[31]),
    .C(_12932_),
    .X(_13087_));
 sky130_fd_sc_hd__inv_2 _23339_ (.A(_13087_),
    .Y(_13088_));
 sky130_fd_sc_hd__nand2_2 _23340_ (.A(_13086_),
    .B(_13088_),
    .Y(_13089_));
 sky130_fd_sc_hd__nand2_2 _23341_ (.A(iY[11]),
    .B(iX[29]),
    .Y(_13090_));
 sky130_fd_sc_hd__xor2_2 _23342_ (.A(_13089_),
    .B(_13090_),
    .X(_13091_));
 sky130_fd_sc_hd__a2bb2o_2 _23343_ (.A1_N(_12933_),
    .A2_N(_12935_),
    .B1(_12602_),
    .B2(_12932_),
    .X(_13093_));
 sky130_fd_sc_hd__xnor2_2 _23344_ (.A(_13091_),
    .B(_13093_),
    .Y(_13094_));
 sky130_fd_sc_hd__nor2_2 _23345_ (.A(_13085_),
    .B(_13094_),
    .Y(_13095_));
 sky130_fd_sc_hd__and2_2 _23346_ (.A(_13085_),
    .B(_13094_),
    .X(_13096_));
 sky130_fd_sc_hd__or2_2 _23347_ (.A(_13095_),
    .B(_13096_),
    .X(_13097_));
 sky130_fd_sc_hd__nor3_2 _23348_ (.A(_12050_),
    .B(_12586_),
    .C(_13097_),
    .Y(_13098_));
 sky130_fd_sc_hd__o21a_2 _23349_ (.A1(_12050_),
    .A2(_12586_),
    .B1(_13097_),
    .X(_13099_));
 sky130_fd_sc_hd__or2_2 _23350_ (.A(_13098_),
    .B(_13099_),
    .X(_13100_));
 sky130_fd_sc_hd__or2b_2 _23351_ (.A(_12937_),
    .B_N(_12936_),
    .X(_13101_));
 sky130_fd_sc_hd__a21bo_2 _23352_ (.A1(_12931_),
    .A2(_12938_),
    .B1_N(_13101_),
    .X(_13102_));
 sky130_fd_sc_hd__xor2_2 _23353_ (.A(_13100_),
    .B(_13102_),
    .X(_13104_));
 sky130_fd_sc_hd__nor2_2 _23354_ (.A(_13076_),
    .B(_13104_),
    .Y(_13105_));
 sky130_fd_sc_hd__and2_2 _23355_ (.A(_13076_),
    .B(_13104_),
    .X(_13106_));
 sky130_fd_sc_hd__nor2_2 _23356_ (.A(_13105_),
    .B(_13106_),
    .Y(_13107_));
 sky130_fd_sc_hd__inv_2 _23357_ (.A(_12980_),
    .Y(_13108_));
 sky130_fd_sc_hd__or2b_2 _23358_ (.A(_12925_),
    .B_N(_12943_),
    .X(_13109_));
 sky130_fd_sc_hd__and4_2 _23359_ (.A(iX[18]),
    .B(iX[19]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_13110_));
 sky130_fd_sc_hd__a22oi_2 _23360_ (.A1(iX[19]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[18]),
    .Y(_13111_));
 sky130_fd_sc_hd__nor2_2 _23361_ (.A(_13110_),
    .B(_13111_),
    .Y(_13112_));
 sky130_fd_sc_hd__nand2_2 _23362_ (.A(iX[17]),
    .B(iY[23]),
    .Y(_13113_));
 sky130_fd_sc_hd__xnor2_2 _23363_ (.A(_13112_),
    .B(_13113_),
    .Y(_13115_));
 sky130_fd_sc_hd__and4_2 _23364_ (.A(iY[18]),
    .B(iY[19]),
    .C(iX[21]),
    .D(iX[22]),
    .X(_13116_));
 sky130_fd_sc_hd__a22oi_2 _23365_ (.A1(iY[19]),
    .A2(iX[21]),
    .B1(iX[22]),
    .B2(iY[18]),
    .Y(_13117_));
 sky130_fd_sc_hd__nor2_2 _23366_ (.A(_13116_),
    .B(_13117_),
    .Y(_13118_));
 sky130_fd_sc_hd__nand2_2 _23367_ (.A(iX[20]),
    .B(iY[20]),
    .Y(_13119_));
 sky130_fd_sc_hd__xnor2_2 _23368_ (.A(_13118_),
    .B(_13119_),
    .Y(_13120_));
 sky130_fd_sc_hd__o21ba_2 _23369_ (.A1(_12957_),
    .A2(_12959_),
    .B1_N(_12956_),
    .X(_13121_));
 sky130_fd_sc_hd__xnor2_2 _23370_ (.A(_13120_),
    .B(_13121_),
    .Y(_13122_));
 sky130_fd_sc_hd__and2_2 _23371_ (.A(_13115_),
    .B(_13122_),
    .X(_13123_));
 sky130_fd_sc_hd__nor2_2 _23372_ (.A(_13115_),
    .B(_13122_),
    .Y(_13124_));
 sky130_fd_sc_hd__or2_2 _23373_ (.A(_13123_),
    .B(_13124_),
    .X(_13126_));
 sky130_fd_sc_hd__or3_2 _23374_ (.A(_12968_),
    .B(_12973_),
    .C(_12974_),
    .X(_13127_));
 sky130_fd_sc_hd__o21ba_2 _23375_ (.A1(_12927_),
    .A2(_12930_),
    .B1_N(_12926_),
    .X(_13128_));
 sky130_fd_sc_hd__and4_2 _23376_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[24]),
    .D(iX[25]),
    .X(_13129_));
 sky130_fd_sc_hd__a22oi_2 _23377_ (.A1(iY[16]),
    .A2(iX[24]),
    .B1(iX[25]),
    .B2(iY[15]),
    .Y(_13130_));
 sky130_fd_sc_hd__nor2_2 _23378_ (.A(_13129_),
    .B(_13130_),
    .Y(_13131_));
 sky130_fd_sc_hd__nand2_2 _23379_ (.A(iY[17]),
    .B(iX[23]),
    .Y(_13132_));
 sky130_fd_sc_hd__xnor2_2 _23380_ (.A(_13131_),
    .B(_13132_),
    .Y(_13133_));
 sky130_fd_sc_hd__xnor2_2 _23381_ (.A(_13128_),
    .B(_13133_),
    .Y(_13134_));
 sky130_fd_sc_hd__o21ai_2 _23382_ (.A1(_12969_),
    .A2(_12974_),
    .B1(_13134_),
    .Y(_13135_));
 sky130_fd_sc_hd__or3_2 _23383_ (.A(_12969_),
    .B(_12974_),
    .C(_13134_),
    .X(_13137_));
 sky130_fd_sc_hd__nand2_2 _23384_ (.A(_13135_),
    .B(_13137_),
    .Y(_13138_));
 sky130_fd_sc_hd__a21oi_2 _23385_ (.A1(_13127_),
    .A2(_12977_),
    .B1(_13138_),
    .Y(_13139_));
 sky130_fd_sc_hd__and3_2 _23386_ (.A(_13127_),
    .B(_12977_),
    .C(_13138_),
    .X(_13140_));
 sky130_fd_sc_hd__or3_2 _23387_ (.A(_13126_),
    .B(_13139_),
    .C(_13140_),
    .X(_13141_));
 sky130_fd_sc_hd__o21ai_2 _23388_ (.A1(_13139_),
    .A2(_13140_),
    .B1(_13126_),
    .Y(_13142_));
 sky130_fd_sc_hd__nand2_2 _23389_ (.A(_13141_),
    .B(_13142_),
    .Y(_13143_));
 sky130_fd_sc_hd__a21oi_2 _23390_ (.A1(_12941_),
    .A2(_13109_),
    .B1(_13143_),
    .Y(_13144_));
 sky130_fd_sc_hd__and3_2 _23391_ (.A(_12941_),
    .B(_13109_),
    .C(_13143_),
    .X(_13145_));
 sky130_fd_sc_hd__a211o_2 _23392_ (.A1(_13108_),
    .A2(_12982_),
    .B1(_13144_),
    .C1(_13145_),
    .X(_13146_));
 sky130_fd_sc_hd__o211ai_2 _23393_ (.A1(_13144_),
    .A2(_13145_),
    .B1(_13108_),
    .C1(_12982_),
    .Y(_13148_));
 sky130_fd_sc_hd__and3_2 _23394_ (.A(_13107_),
    .B(_13146_),
    .C(_13148_),
    .X(_13149_));
 sky130_fd_sc_hd__a21oi_2 _23395_ (.A1(_13146_),
    .A2(_13148_),
    .B1(_13107_),
    .Y(_13150_));
 sky130_fd_sc_hd__a211o_2 _23396_ (.A1(_13075_),
    .A2(_12990_),
    .B1(_13149_),
    .C1(_13150_),
    .X(_13151_));
 sky130_fd_sc_hd__o211ai_2 _23397_ (.A1(_13149_),
    .A2(_13150_),
    .B1(_13075_),
    .C1(_12990_),
    .Y(_13152_));
 sky130_fd_sc_hd__inv_2 _23398_ (.A(_13036_),
    .Y(_13153_));
 sky130_fd_sc_hd__or2b_2 _23399_ (.A(_12986_),
    .B_N(_12988_),
    .X(_13154_));
 sky130_fd_sc_hd__inv_2 _23400_ (.A(_13154_),
    .Y(_13155_));
 sky130_fd_sc_hd__and4_2 _23401_ (.A(iX[12]),
    .B(iX[13]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_13156_));
 sky130_fd_sc_hd__a22oi_2 _23402_ (.A1(iX[13]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[12]),
    .Y(_13157_));
 sky130_fd_sc_hd__nor2_2 _23403_ (.A(_13156_),
    .B(_13157_),
    .Y(_13159_));
 sky130_fd_sc_hd__nand2_2 _23404_ (.A(iX[11]),
    .B(iY[29]),
    .Y(_13160_));
 sky130_fd_sc_hd__xnor2_2 _23405_ (.A(_13159_),
    .B(_13160_),
    .Y(_13161_));
 sky130_fd_sc_hd__o21ba_2 _23406_ (.A1(_12999_),
    .A2(_13001_),
    .B1_N(_12998_),
    .X(_13162_));
 sky130_fd_sc_hd__xnor2_2 _23407_ (.A(_13161_),
    .B(_13162_),
    .Y(_13163_));
 sky130_fd_sc_hd__nand3_2 _23408_ (.A(iX[10]),
    .B(iY[30]),
    .C(_13163_),
    .Y(_13164_));
 sky130_fd_sc_hd__a21o_2 _23409_ (.A1(iX[10]),
    .A2(iY[30]),
    .B1(_13163_),
    .X(_13165_));
 sky130_fd_sc_hd__nand2_2 _23410_ (.A(_13164_),
    .B(_13165_),
    .Y(_13166_));
 sky130_fd_sc_hd__or2b_2 _23411_ (.A(_13003_),
    .B_N(_13002_),
    .X(_13167_));
 sky130_fd_sc_hd__nand2_2 _23412_ (.A(_13167_),
    .B(_13008_),
    .Y(_13168_));
 sky130_fd_sc_hd__xnor2_2 _23413_ (.A(_13166_),
    .B(_13168_),
    .Y(_13170_));
 sky130_fd_sc_hd__and2_2 _23414_ (.A(iX[9]),
    .B(iY[31]),
    .X(_13171_));
 sky130_fd_sc_hd__nor2_2 _23415_ (.A(_13170_),
    .B(_13171_),
    .Y(_13172_));
 sky130_fd_sc_hd__and2_2 _23416_ (.A(_13170_),
    .B(_13171_),
    .X(_13173_));
 sky130_fd_sc_hd__nor2_2 _23417_ (.A(_13172_),
    .B(_13173_),
    .Y(_13174_));
 sky130_fd_sc_hd__or2b_2 _23418_ (.A(_13020_),
    .B_N(_13025_),
    .X(_13175_));
 sky130_fd_sc_hd__or2b_2 _23419_ (.A(_13019_),
    .B_N(_13026_),
    .X(_13176_));
 sky130_fd_sc_hd__and2b_2 _23420_ (.A_N(_12962_),
    .B(_12960_),
    .X(_13177_));
 sky130_fd_sc_hd__o21ba_2 _23421_ (.A1(_13022_),
    .A2(_13024_),
    .B1_N(_13021_),
    .X(_13178_));
 sky130_fd_sc_hd__o21ba_2 _23422_ (.A1(_12952_),
    .A2(_12954_),
    .B1_N(_12951_),
    .X(_13179_));
 sky130_fd_sc_hd__and4_2 _23423_ (.A(iX[15]),
    .B(iX[16]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_13181_));
 sky130_fd_sc_hd__a22oi_2 _23424_ (.A1(iX[16]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[15]),
    .Y(_13182_));
 sky130_fd_sc_hd__nor2_2 _23425_ (.A(_13181_),
    .B(_13182_),
    .Y(_13183_));
 sky130_fd_sc_hd__nand2_2 _23426_ (.A(iX[14]),
    .B(iY[26]),
    .Y(_13184_));
 sky130_fd_sc_hd__xnor2_2 _23427_ (.A(_13183_),
    .B(_13184_),
    .Y(_13185_));
 sky130_fd_sc_hd__xnor2_2 _23428_ (.A(_13179_),
    .B(_13185_),
    .Y(_13186_));
 sky130_fd_sc_hd__xnor2_2 _23429_ (.A(_13178_),
    .B(_13186_),
    .Y(_13187_));
 sky130_fd_sc_hd__o21a_2 _23430_ (.A1(_13177_),
    .A2(_12964_),
    .B1(_13187_),
    .X(_13188_));
 sky130_fd_sc_hd__nor3_2 _23431_ (.A(_13177_),
    .B(_12964_),
    .C(_13187_),
    .Y(_13189_));
 sky130_fd_sc_hd__a211oi_2 _23432_ (.A1(_13175_),
    .A2(_13176_),
    .B1(_13188_),
    .C1(_13189_),
    .Y(_13190_));
 sky130_fd_sc_hd__o211a_2 _23433_ (.A1(_13188_),
    .A2(_13189_),
    .B1(_13175_),
    .C1(_13176_),
    .X(_13192_));
 sky130_fd_sc_hd__nor2_2 _23434_ (.A(_13029_),
    .B(_13031_),
    .Y(_13193_));
 sky130_fd_sc_hd__or3_2 _23435_ (.A(_13190_),
    .B(_13192_),
    .C(_13193_),
    .X(_13194_));
 sky130_fd_sc_hd__o21ai_2 _23436_ (.A1(_13190_),
    .A2(_13192_),
    .B1(_13193_),
    .Y(_13195_));
 sky130_fd_sc_hd__and3_2 _23437_ (.A(_13174_),
    .B(_13194_),
    .C(_13195_),
    .X(_13196_));
 sky130_fd_sc_hd__a21oi_2 _23438_ (.A1(_13194_),
    .A2(_13195_),
    .B1(_13174_),
    .Y(_13197_));
 sky130_fd_sc_hd__or3_2 _23439_ (.A(_13155_),
    .B(_13196_),
    .C(_13197_),
    .X(_13198_));
 sky130_fd_sc_hd__o21ai_2 _23440_ (.A1(_13196_),
    .A2(_13197_),
    .B1(_13155_),
    .Y(_13199_));
 sky130_fd_sc_hd__nand2_2 _23441_ (.A(_13198_),
    .B(_13199_),
    .Y(_13200_));
 sky130_fd_sc_hd__a21o_2 _23442_ (.A1(_13034_),
    .A2(_13153_),
    .B1(_13200_),
    .X(_13201_));
 sky130_fd_sc_hd__nand3_2 _23443_ (.A(_13034_),
    .B(_13153_),
    .C(_13200_),
    .Y(_13203_));
 sky130_fd_sc_hd__nand4_2 _23444_ (.A(_13151_),
    .B(_13152_),
    .C(_13201_),
    .D(_13203_),
    .Y(_13204_));
 sky130_fd_sc_hd__a22o_2 _23445_ (.A1(_13151_),
    .A2(_13152_),
    .B1(_13201_),
    .B2(_13203_),
    .X(_13205_));
 sky130_fd_sc_hd__o211a_2 _23446_ (.A1(_12993_),
    .A2(_13074_),
    .B1(_13204_),
    .C1(_13205_),
    .X(_13206_));
 sky130_fd_sc_hd__a211oi_2 _23447_ (.A1(_13204_),
    .A2(_13205_),
    .B1(_12993_),
    .C1(_13074_),
    .Y(_13207_));
 sky130_fd_sc_hd__or2_2 _23448_ (.A(_13206_),
    .B(_13207_),
    .X(_13208_));
 sky130_fd_sc_hd__nand2_2 _23449_ (.A(_13040_),
    .B(_13042_),
    .Y(_13209_));
 sky130_fd_sc_hd__xnor2_2 _23450_ (.A(_13208_),
    .B(_13209_),
    .Y(_13210_));
 sky130_fd_sc_hd__o21a_2 _23451_ (.A1(_13047_),
    .A2(_13050_),
    .B1(_13210_),
    .X(_13211_));
 sky130_fd_sc_hd__nor3_2 _23452_ (.A(_13047_),
    .B(_13050_),
    .C(_13210_),
    .Y(_13212_));
 sky130_fd_sc_hd__nor2_2 _23453_ (.A(_13211_),
    .B(_13212_),
    .Y(_13214_));
 sky130_fd_sc_hd__a31o_2 _23454_ (.A1(iX[8]),
    .A2(iY[31]),
    .A3(_13012_),
    .B1(_13010_),
    .X(_13215_));
 sky130_fd_sc_hd__xnor2_2 _23455_ (.A(_13214_),
    .B(_13215_),
    .Y(_13216_));
 sky130_fd_sc_hd__nor2_2 _23456_ (.A(_13053_),
    .B(_13055_),
    .Y(_13217_));
 sky130_fd_sc_hd__or2_2 _23457_ (.A(_13216_),
    .B(_13217_),
    .X(_13218_));
 sky130_fd_sc_hd__nand2_2 _23458_ (.A(_13216_),
    .B(_13217_),
    .Y(_13219_));
 sky130_fd_sc_hd__nand2_2 _23459_ (.A(_13218_),
    .B(_13219_),
    .Y(_13220_));
 sky130_fd_sc_hd__or2_2 _23460_ (.A(_12200_),
    .B(_12442_),
    .X(_13221_));
 sky130_fd_sc_hd__or4b_2 _23461_ (.A(_12443_),
    .B(_12693_),
    .C(_13061_),
    .D_N(_13221_),
    .X(_13222_));
 sky130_fd_sc_hd__or2b_2 _23462_ (.A(_13058_),
    .B_N(_12691_),
    .X(_13223_));
 sky130_fd_sc_hd__and3b_2 _23463_ (.A_N(_13059_),
    .B(_13222_),
    .C(_13223_),
    .X(_13225_));
 sky130_fd_sc_hd__nand2_2 _23464_ (.A(_12445_),
    .B(_12444_),
    .Y(_13226_));
 sky130_fd_sc_hd__o31a_2 _23465_ (.A1(_12693_),
    .A2(_13061_),
    .A3(_13226_),
    .B1(_13225_),
    .X(_13227_));
 sky130_fd_sc_hd__a31oi_2 _23466_ (.A1(_12204_),
    .A2(_12209_),
    .A3(_13225_),
    .B1(_13227_),
    .Y(_13228_));
 sky130_fd_sc_hd__xor2_2 _23467_ (.A(_13220_),
    .B(_13228_),
    .X(_13229_));
 sky130_fd_sc_hd__or2b_2 _23468_ (.A(_12854_),
    .B_N(_12839_),
    .X(_13230_));
 sky130_fd_sc_hd__or2_2 _23469_ (.A(_12746_),
    .B(_12747_),
    .X(_13231_));
 sky130_fd_sc_hd__and4_2 _23470_ (.A(_12217_),
    .B(_12454_),
    .C(_12742_),
    .D(_12805_),
    .X(_13232_));
 sky130_fd_sc_hd__o211a_2 _23471_ (.A1(iX[7]),
    .A2(iX[39]),
    .B1(iX[38]),
    .C1(iX[6]),
    .X(_13233_));
 sky130_fd_sc_hd__a21o_2 _23472_ (.A1(iX[7]),
    .A2(iX[39]),
    .B1(_13233_),
    .X(_13234_));
 sky130_fd_sc_hd__a41o_2 _23473_ (.A1(_12453_),
    .A2(_12742_),
    .A3(_12744_),
    .A4(_12805_),
    .B1(_13234_),
    .X(_13236_));
 sky130_fd_sc_hd__a21o_4 _23474_ (.A1(_12222_),
    .A2(_13232_),
    .B1(_13236_),
    .X(_13237_));
 sky130_fd_sc_hd__and2_2 _23475_ (.A(iX[8]),
    .B(iX[40]),
    .X(_13238_));
 sky130_fd_sc_hd__nor2_2 _23476_ (.A(iX[8]),
    .B(iX[40]),
    .Y(_13239_));
 sky130_fd_sc_hd__nor2_2 _23477_ (.A(_13238_),
    .B(_13239_),
    .Y(_13240_));
 sky130_fd_sc_hd__xnor2_2 _23478_ (.A(_13237_),
    .B(_13240_),
    .Y(_13241_));
 sky130_fd_sc_hd__nor2_2 _23479_ (.A(_11574_),
    .B(_13241_),
    .Y(_13242_));
 sky130_fd_sc_hd__and3_2 _23480_ (.A(_11378_),
    .B(_12811_),
    .C(_13242_),
    .X(_13243_));
 sky130_fd_sc_hd__xor2_2 _23481_ (.A(_13237_),
    .B(_13240_),
    .X(_13244_));
 sky130_fd_sc_hd__a22o_2 _23482_ (.A1(_11582_),
    .A2(_12811_),
    .B1(_13244_),
    .B2(_11378_),
    .X(_13245_));
 sky130_fd_sc_hd__or4b_4 _23483_ (.A(_11791_),
    .B(_13231_),
    .C(_13243_),
    .D_N(_13245_),
    .X(_13247_));
 sky130_fd_sc_hd__or3b_2 _23484_ (.A(_11565_),
    .B(_12808_),
    .C_N(_13242_),
    .X(_13248_));
 sky130_fd_sc_hd__a22o_2 _23485_ (.A1(_12450_),
    .A2(_12810_),
    .B1(_13248_),
    .B2(_13245_),
    .X(_13249_));
 sky130_fd_sc_hd__a31o_2 _23486_ (.A1(_12450_),
    .A2(_12460_),
    .A3(_12812_),
    .B1(_12809_),
    .X(_13250_));
 sky130_fd_sc_hd__nand3_2 _23487_ (.A(_13247_),
    .B(_13249_),
    .C(_13250_),
    .Y(_13251_));
 sky130_fd_sc_hd__a21o_2 _23488_ (.A1(_13247_),
    .A2(_13249_),
    .B1(_13250_),
    .X(_13252_));
 sky130_fd_sc_hd__nor2_2 _23489_ (.A(_12244_),
    .B(_12456_),
    .Y(_13253_));
 sky130_fd_sc_hd__xnor2_2 _23490_ (.A(_12823_),
    .B(_13253_),
    .Y(_13254_));
 sky130_fd_sc_hd__nand2_2 _23491_ (.A(_11829_),
    .B(_12477_),
    .Y(_13255_));
 sky130_fd_sc_hd__xnor2_2 _23492_ (.A(_13254_),
    .B(_13255_),
    .Y(_13256_));
 sky130_fd_sc_hd__nand3_2 _23493_ (.A(_13251_),
    .B(_13252_),
    .C(_13256_),
    .Y(_13258_));
 sky130_fd_sc_hd__a21o_2 _23494_ (.A1(_13251_),
    .A2(_13252_),
    .B1(_13256_),
    .X(_13259_));
 sky130_fd_sc_hd__a21bo_2 _23495_ (.A1(_12821_),
    .A2(_12830_),
    .B1_N(_12820_),
    .X(_13260_));
 sky130_fd_sc_hd__nand3_2 _23496_ (.A(_13258_),
    .B(_13259_),
    .C(_13260_),
    .Y(_13261_));
 sky130_fd_sc_hd__a21o_2 _23497_ (.A1(_13258_),
    .A2(_13259_),
    .B1(_13260_),
    .X(_13262_));
 sky130_fd_sc_hd__a31o_2 _23498_ (.A1(_12827_),
    .A2(_12759_),
    .A3(_12826_),
    .B1(_12824_),
    .X(_13263_));
 sky130_fd_sc_hd__nor2_2 _23499_ (.A(_12227_),
    .B(_12772_),
    .Y(_13264_));
 sky130_fd_sc_hd__or3b_2 _23500_ (.A(_11569_),
    .B(_12849_),
    .C_N(_13264_),
    .X(_13265_));
 sky130_fd_sc_hd__a21o_2 _23501_ (.A1(_11581_),
    .A2(_12845_),
    .B1(_13264_),
    .X(_13266_));
 sky130_fd_sc_hd__xor2_2 _23502_ (.A(iY[8]),
    .B(iY[40]),
    .X(_13267_));
 sky130_fd_sc_hd__a21boi_2 _23503_ (.A1(_12767_),
    .A2(_12841_),
    .B1_N(_12842_),
    .Y(_13269_));
 sky130_fd_sc_hd__and2_2 _23504_ (.A(iY[7]),
    .B(iY[39]),
    .X(_13270_));
 sky130_fd_sc_hd__o21a_2 _23505_ (.A1(_12768_),
    .A2(_13270_),
    .B1(_12842_),
    .X(_13271_));
 sky130_fd_sc_hd__o21a_2 _23506_ (.A1(_12771_),
    .A2(_13269_),
    .B1(_13271_),
    .X(_13272_));
 sky130_fd_sc_hd__xnor2_2 _23507_ (.A(_13267_),
    .B(_13272_),
    .Y(_13273_));
 sky130_fd_sc_hd__inv_2 _23508_ (.A(_13273_),
    .Y(_13274_));
 sky130_fd_sc_hd__nand4_2 _23509_ (.A(_11373_),
    .B(_13265_),
    .C(_13266_),
    .D(_13274_),
    .Y(_13275_));
 sky130_fd_sc_hd__a22o_2 _23510_ (.A1(_13265_),
    .A2(_13266_),
    .B1(_13274_),
    .B2(_11374_),
    .X(_13276_));
 sky130_fd_sc_hd__nand3_2 _23511_ (.A(_13263_),
    .B(_13275_),
    .C(_13276_),
    .Y(_13277_));
 sky130_fd_sc_hd__a21o_2 _23512_ (.A1(_13275_),
    .A2(_13276_),
    .B1(_13263_),
    .X(_13278_));
 sky130_fd_sc_hd__a21o_2 _23513_ (.A1(_13277_),
    .A2(_13278_),
    .B1(_12847_),
    .X(_13280_));
 sky130_fd_sc_hd__nand3_2 _23514_ (.A(_12847_),
    .B(_13277_),
    .C(_13278_),
    .Y(_13281_));
 sky130_fd_sc_hd__nand4_2 _23515_ (.A(_13261_),
    .B(_13262_),
    .C(_13280_),
    .D(_13281_),
    .Y(_13282_));
 sky130_fd_sc_hd__a22o_2 _23516_ (.A1(_13261_),
    .A2(_13262_),
    .B1(_13280_),
    .B2(_13281_),
    .X(_13283_));
 sky130_fd_sc_hd__o211a_2 _23517_ (.A1(_12836_),
    .A2(_12856_),
    .B1(_13282_),
    .C1(_13283_),
    .X(_13284_));
 sky130_fd_sc_hd__a211oi_2 _23518_ (.A1(_13282_),
    .A2(_13283_),
    .B1(_12836_),
    .C1(_12856_),
    .Y(_13285_));
 sky130_fd_sc_hd__nor3_2 _23519_ (.A(_13230_),
    .B(_13284_),
    .C(_13285_),
    .Y(_13286_));
 sky130_fd_sc_hd__o21a_2 _23520_ (.A1(_13284_),
    .A2(_13285_),
    .B1(_13230_),
    .X(_13287_));
 sky130_fd_sc_hd__nor2_2 _23521_ (.A(_13286_),
    .B(_13287_),
    .Y(_13288_));
 sky130_fd_sc_hd__nand2_2 _23522_ (.A(_12858_),
    .B(_12860_),
    .Y(_13289_));
 sky130_fd_sc_hd__xor2_2 _23523_ (.A(_13288_),
    .B(_13289_),
    .X(_13291_));
 sky130_fd_sc_hd__o21ba_2 _23524_ (.A1(_12784_),
    .A2(_12864_),
    .B1_N(_12863_),
    .X(_13292_));
 sky130_fd_sc_hd__xnor2_2 _23525_ (.A(_13291_),
    .B(_13292_),
    .Y(_13293_));
 sky130_fd_sc_hd__or2_2 _23526_ (.A(_12863_),
    .B(_12864_),
    .X(_13294_));
 sky130_fd_sc_hd__nor2_2 _23527_ (.A(_12783_),
    .B(_13294_),
    .Y(_13295_));
 sky130_fd_sc_hd__xnor2_2 _23528_ (.A(_13293_),
    .B(_13295_),
    .Y(_13296_));
 sky130_fd_sc_hd__nor2_2 _23529_ (.A(_12733_),
    .B(_12904_),
    .Y(_13297_));
 sky130_fd_sc_hd__and4_2 _23530_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[37]),
    .D(iX[38]),
    .X(_13298_));
 sky130_fd_sc_hd__a22oi_2 _23531_ (.A1(iY[35]),
    .A2(iX[37]),
    .B1(iX[38]),
    .B2(iY[34]),
    .Y(_13299_));
 sky130_fd_sc_hd__nand2_2 _23532_ (.A(iY[33]),
    .B(iX[39]),
    .Y(_13300_));
 sky130_fd_sc_hd__or3_2 _23533_ (.A(_13298_),
    .B(_13299_),
    .C(_13300_),
    .X(_13302_));
 sky130_fd_sc_hd__o21ai_2 _23534_ (.A1(_13298_),
    .A2(_13299_),
    .B1(_13300_),
    .Y(_13303_));
 sky130_fd_sc_hd__o21bai_2 _23535_ (.A1(_12869_),
    .A2(_12870_),
    .B1_N(_12868_),
    .Y(_13304_));
 sky130_fd_sc_hd__nand3_2 _23536_ (.A(_13302_),
    .B(_13303_),
    .C(_13304_),
    .Y(_13305_));
 sky130_fd_sc_hd__a21o_2 _23537_ (.A1(_13302_),
    .A2(_13303_),
    .B1(_13304_),
    .X(_13306_));
 sky130_fd_sc_hd__and4_2 _23538_ (.A(iY[32]),
    .B(iX[36]),
    .C(iY[36]),
    .D(iX[40]),
    .X(_13307_));
 sky130_fd_sc_hd__a22oi_2 _23539_ (.A1(iX[36]),
    .A2(iY[36]),
    .B1(iX[40]),
    .B2(iY[32]),
    .Y(_13308_));
 sky130_fd_sc_hd__nor2_2 _23540_ (.A(_13307_),
    .B(_13308_),
    .Y(_13309_));
 sky130_fd_sc_hd__nand2_2 _23541_ (.A(iX[35]),
    .B(iY[37]),
    .Y(_13310_));
 sky130_fd_sc_hd__xnor2_2 _23542_ (.A(_13309_),
    .B(_13310_),
    .Y(_13311_));
 sky130_fd_sc_hd__nand3_2 _23543_ (.A(_13305_),
    .B(_13306_),
    .C(_13311_),
    .Y(_13313_));
 sky130_fd_sc_hd__a21o_2 _23544_ (.A1(_13305_),
    .A2(_13306_),
    .B1(_13311_),
    .X(_13314_));
 sky130_fd_sc_hd__a21bo_2 _23545_ (.A1(_12876_),
    .A2(_12881_),
    .B1_N(_12875_),
    .X(_13315_));
 sky130_fd_sc_hd__and3_2 _23546_ (.A(_13313_),
    .B(_13314_),
    .C(_13315_),
    .X(_13316_));
 sky130_fd_sc_hd__a21oi_2 _23547_ (.A1(_13313_),
    .A2(_13314_),
    .B1(_13315_),
    .Y(_13317_));
 sky130_fd_sc_hd__a31o_2 _23548_ (.A1(iX[34]),
    .A2(iY[37]),
    .A3(_12878_),
    .B1(_12877_),
    .X(_13318_));
 sky130_fd_sc_hd__and4_2 _23549_ (.A(iX[33]),
    .B(iX[34]),
    .C(iY[38]),
    .D(iY[39]),
    .X(_13319_));
 sky130_fd_sc_hd__a22oi_2 _23550_ (.A1(iX[34]),
    .A2(iY[38]),
    .B1(iY[39]),
    .B2(iX[33]),
    .Y(_13320_));
 sky130_fd_sc_hd__nor2_2 _23551_ (.A(_13319_),
    .B(_13320_),
    .Y(_13321_));
 sky130_fd_sc_hd__nand2_2 _23552_ (.A(iX[32]),
    .B(iY[40]),
    .Y(_13322_));
 sky130_fd_sc_hd__xnor2_2 _23553_ (.A(_13321_),
    .B(_13322_),
    .Y(_13324_));
 sky130_fd_sc_hd__xor2_2 _23554_ (.A(_13318_),
    .B(_13324_),
    .X(_13325_));
 sky130_fd_sc_hd__xnor2_2 _23555_ (.A(_12888_),
    .B(_13325_),
    .Y(_13326_));
 sky130_fd_sc_hd__nor3_2 _23556_ (.A(_13316_),
    .B(_13317_),
    .C(_13326_),
    .Y(_13327_));
 sky130_fd_sc_hd__o21a_2 _23557_ (.A1(_13316_),
    .A2(_13317_),
    .B1(_13326_),
    .X(_13328_));
 sky130_fd_sc_hd__a211oi_2 _23558_ (.A1(_12886_),
    .A2(_12896_),
    .B1(_13327_),
    .C1(_13328_),
    .Y(_13329_));
 sky130_fd_sc_hd__o211a_2 _23559_ (.A1(_13327_),
    .A2(_13328_),
    .B1(_12886_),
    .C1(_12896_),
    .X(_13330_));
 sky130_fd_sc_hd__o21ba_2 _23560_ (.A1(_13329_),
    .A2(_13330_),
    .B1_N(_12892_),
    .X(_13331_));
 sky130_fd_sc_hd__nor3b_2 _23561_ (.A(_13329_),
    .B(_13330_),
    .C_N(_12892_),
    .Y(_13332_));
 sky130_fd_sc_hd__nor2_2 _23562_ (.A(_13331_),
    .B(_13332_),
    .Y(_13333_));
 sky130_fd_sc_hd__nand2_2 _23563_ (.A(_12898_),
    .B(_12900_),
    .Y(_13334_));
 sky130_fd_sc_hd__xnor2_2 _23564_ (.A(_13333_),
    .B(_13334_),
    .Y(_13335_));
 sky130_fd_sc_hd__a21bo_2 _23565_ (.A1(_12729_),
    .A2(_12903_),
    .B1_N(_12902_),
    .X(_13336_));
 sky130_fd_sc_hd__xor2_2 _23566_ (.A(_13335_),
    .B(_13336_),
    .X(_13337_));
 sky130_fd_sc_hd__xnor2_2 _23567_ (.A(_13297_),
    .B(_13337_),
    .Y(_13338_));
 sky130_fd_sc_hd__and3b_2 _23568_ (.A_N(_12908_),
    .B(_13338_),
    .C(_12736_),
    .X(_13339_));
 sky130_fd_sc_hd__nor2_2 _23569_ (.A(_12909_),
    .B(_13338_),
    .Y(_13340_));
 sky130_fd_sc_hd__nor2_2 _23570_ (.A(_13339_),
    .B(_13340_),
    .Y(_13341_));
 sky130_fd_sc_hd__xnor2_2 _23571_ (.A(_13296_),
    .B(_13341_),
    .Y(_13342_));
 sky130_fd_sc_hd__xnor2_2 _23572_ (.A(oO[8]),
    .B(_13342_),
    .Y(_13343_));
 sky130_fd_sc_hd__a21boi_2 _23573_ (.A1(_12327_),
    .A2(_12913_),
    .B1_N(_12912_),
    .Y(_13345_));
 sky130_fd_sc_hd__xnor2_2 _23574_ (.A(_13343_),
    .B(_13345_),
    .Y(_13346_));
 sky130_fd_sc_hd__nand2_2 _23575_ (.A(_12915_),
    .B(_12918_),
    .Y(_13347_));
 sky130_fd_sc_hd__o21ai_2 _23576_ (.A1(_12919_),
    .A2(_12921_),
    .B1(_13347_),
    .Y(_13348_));
 sky130_fd_sc_hd__xnor2_2 _23577_ (.A(_13346_),
    .B(_13348_),
    .Y(_13349_));
 sky130_fd_sc_hd__xnor2_2 _23578_ (.A(_13229_),
    .B(_13349_),
    .Y(_13350_));
 sky130_fd_sc_hd__xor2_2 _23579_ (.A(_13073_),
    .B(_13350_),
    .X(oO[40]));
 sky130_fd_sc_hd__and2b_2 _23580_ (.A_N(_13208_),
    .B(_13209_),
    .X(_13351_));
 sky130_fd_sc_hd__and2_2 _23581_ (.A(_13091_),
    .B(_13093_),
    .X(_13352_));
 sky130_fd_sc_hd__and3_2 _23582_ (.A(iY[11]),
    .B(iX[31]),
    .C(_12932_),
    .X(_13353_));
 sky130_fd_sc_hd__a22oi_2 _23583_ (.A1(iY[11]),
    .A2(iX[30]),
    .B1(iX[31]),
    .B2(iY[10]),
    .Y(_13355_));
 sky130_fd_sc_hd__or2_2 _23584_ (.A(_13353_),
    .B(_13355_),
    .X(_13356_));
 sky130_fd_sc_hd__a31o_2 _23585_ (.A1(iY[11]),
    .A2(iX[29]),
    .A3(_13086_),
    .B1(_13087_),
    .X(_13357_));
 sky130_fd_sc_hd__xnor2_2 _23586_ (.A(_13356_),
    .B(_13357_),
    .Y(_13358_));
 sky130_fd_sc_hd__and4_2 _23587_ (.A(iY[12]),
    .B(iY[13]),
    .C(iX[28]),
    .D(iX[29]),
    .X(_13359_));
 sky130_fd_sc_hd__a22oi_2 _23588_ (.A1(iY[13]),
    .A2(iX[28]),
    .B1(iX[29]),
    .B2(iY[12]),
    .Y(_13360_));
 sky130_fd_sc_hd__nor2_2 _23589_ (.A(_13359_),
    .B(_13360_),
    .Y(_13361_));
 sky130_fd_sc_hd__nand2_2 _23590_ (.A(iY[14]),
    .B(iX[27]),
    .Y(_13362_));
 sky130_fd_sc_hd__xnor2_2 _23591_ (.A(_13361_),
    .B(_13362_),
    .Y(_13363_));
 sky130_fd_sc_hd__nand2_2 _23592_ (.A(_13358_),
    .B(_13363_),
    .Y(_13364_));
 sky130_fd_sc_hd__or2_2 _23593_ (.A(_13358_),
    .B(_13363_),
    .X(_13366_));
 sky130_fd_sc_hd__and2_2 _23594_ (.A(_13364_),
    .B(_13366_),
    .X(_13367_));
 sky130_fd_sc_hd__o21a_2 _23595_ (.A1(_13352_),
    .A2(_13095_),
    .B1(_13367_),
    .X(_13368_));
 sky130_fd_sc_hd__nor3_2 _23596_ (.A(_13352_),
    .B(_13095_),
    .C(_13367_),
    .Y(_13369_));
 sky130_fd_sc_hd__or2_2 _23597_ (.A(_13368_),
    .B(_13369_),
    .X(_13370_));
 sky130_fd_sc_hd__inv_2 _23598_ (.A(_13139_),
    .Y(_13371_));
 sky130_fd_sc_hd__and2b_2 _23599_ (.A_N(_13100_),
    .B(_13102_),
    .X(_13372_));
 sky130_fd_sc_hd__and4_2 _23600_ (.A(iX[19]),
    .B(iX[20]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_13373_));
 sky130_fd_sc_hd__a22oi_2 _23601_ (.A1(iX[20]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[19]),
    .Y(_13374_));
 sky130_fd_sc_hd__nor2_2 _23602_ (.A(_13373_),
    .B(_13374_),
    .Y(_13375_));
 sky130_fd_sc_hd__nand2_2 _23603_ (.A(iX[18]),
    .B(iY[23]),
    .Y(_13377_));
 sky130_fd_sc_hd__xnor2_2 _23604_ (.A(_13375_),
    .B(_13377_),
    .Y(_13378_));
 sky130_fd_sc_hd__and4_2 _23605_ (.A(iY[18]),
    .B(iY[19]),
    .C(iX[22]),
    .D(iX[23]),
    .X(_13379_));
 sky130_fd_sc_hd__a22oi_2 _23606_ (.A1(iY[19]),
    .A2(iX[22]),
    .B1(iX[23]),
    .B2(iY[18]),
    .Y(_13380_));
 sky130_fd_sc_hd__nor2_2 _23607_ (.A(_13379_),
    .B(_13380_),
    .Y(_13381_));
 sky130_fd_sc_hd__nand2_2 _23608_ (.A(iY[20]),
    .B(iX[21]),
    .Y(_13382_));
 sky130_fd_sc_hd__xnor2_2 _23609_ (.A(_13381_),
    .B(_13382_),
    .Y(_13383_));
 sky130_fd_sc_hd__o21ba_2 _23610_ (.A1(_13117_),
    .A2(_13119_),
    .B1_N(_13116_),
    .X(_13384_));
 sky130_fd_sc_hd__xnor2_2 _23611_ (.A(_13383_),
    .B(_13384_),
    .Y(_13385_));
 sky130_fd_sc_hd__and2_2 _23612_ (.A(_13378_),
    .B(_13385_),
    .X(_13386_));
 sky130_fd_sc_hd__nor2_2 _23613_ (.A(_13378_),
    .B(_13385_),
    .Y(_13388_));
 sky130_fd_sc_hd__or2_2 _23614_ (.A(_13386_),
    .B(_13388_),
    .X(_13389_));
 sky130_fd_sc_hd__or2b_2 _23615_ (.A(_13128_),
    .B_N(_13133_),
    .X(_13390_));
 sky130_fd_sc_hd__a31o_2 _23616_ (.A1(iY[17]),
    .A2(iX[23]),
    .A3(_13131_),
    .B1(_13129_),
    .X(_13391_));
 sky130_fd_sc_hd__and4_2 _23617_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[25]),
    .D(iX[26]),
    .X(_13392_));
 sky130_fd_sc_hd__a22oi_2 _23618_ (.A1(iY[16]),
    .A2(iX[25]),
    .B1(iX[26]),
    .B2(iY[15]),
    .Y(_13393_));
 sky130_fd_sc_hd__and4bb_2 _23619_ (.A_N(_13392_),
    .B_N(_13393_),
    .C(iY[17]),
    .D(iX[24]),
    .X(_13394_));
 sky130_fd_sc_hd__o2bb2a_2 _23620_ (.A1_N(iY[17]),
    .A2_N(iX[24]),
    .B1(_13392_),
    .B2(_13393_),
    .X(_13395_));
 sky130_fd_sc_hd__nor2_2 _23621_ (.A(_13394_),
    .B(_13395_),
    .Y(_13396_));
 sky130_fd_sc_hd__o21ai_2 _23622_ (.A1(_13077_),
    .A2(_13082_),
    .B1(_13396_),
    .Y(_13397_));
 sky130_fd_sc_hd__or3_2 _23623_ (.A(_13077_),
    .B(_13082_),
    .C(_13396_),
    .X(_13399_));
 sky130_fd_sc_hd__and2_2 _23624_ (.A(_13397_),
    .B(_13399_),
    .X(_13400_));
 sky130_fd_sc_hd__xnor2_2 _23625_ (.A(_13391_),
    .B(_13400_),
    .Y(_13401_));
 sky130_fd_sc_hd__a21oi_2 _23626_ (.A1(_13390_),
    .A2(_13135_),
    .B1(_13401_),
    .Y(_13402_));
 sky130_fd_sc_hd__and3_2 _23627_ (.A(_13390_),
    .B(_13135_),
    .C(_13401_),
    .X(_13403_));
 sky130_fd_sc_hd__or3_2 _23628_ (.A(_13389_),
    .B(_13402_),
    .C(_13403_),
    .X(_13404_));
 sky130_fd_sc_hd__o21ai_2 _23629_ (.A1(_13402_),
    .A2(_13403_),
    .B1(_13389_),
    .Y(_13405_));
 sky130_fd_sc_hd__o211a_2 _23630_ (.A1(_13098_),
    .A2(_13372_),
    .B1(_13404_),
    .C1(_13405_),
    .X(_13406_));
 sky130_fd_sc_hd__a211oi_2 _23631_ (.A1(_13404_),
    .A2(_13405_),
    .B1(_13098_),
    .C1(_13372_),
    .Y(_13407_));
 sky130_fd_sc_hd__a211oi_2 _23632_ (.A1(_13371_),
    .A2(_13141_),
    .B1(_13406_),
    .C1(_13407_),
    .Y(_13408_));
 sky130_fd_sc_hd__o211a_2 _23633_ (.A1(_13406_),
    .A2(_13407_),
    .B1(_13371_),
    .C1(_13141_),
    .X(_13410_));
 sky130_fd_sc_hd__or3_2 _23634_ (.A(_13370_),
    .B(_13408_),
    .C(_13410_),
    .X(_13411_));
 sky130_fd_sc_hd__o21ai_2 _23635_ (.A1(_13408_),
    .A2(_13410_),
    .B1(_13370_),
    .Y(_13412_));
 sky130_fd_sc_hd__o211ai_2 _23636_ (.A1(_13105_),
    .A2(_13149_),
    .B1(_13411_),
    .C1(_13412_),
    .Y(_13413_));
 sky130_fd_sc_hd__a211o_2 _23637_ (.A1(_13411_),
    .A2(_13412_),
    .B1(_13105_),
    .C1(_13149_),
    .X(_13414_));
 sky130_fd_sc_hd__inv_2 _23638_ (.A(_13196_),
    .Y(_13415_));
 sky130_fd_sc_hd__or2b_2 _23639_ (.A(_13144_),
    .B_N(_13146_),
    .X(_13416_));
 sky130_fd_sc_hd__inv_2 _23640_ (.A(_13416_),
    .Y(_13417_));
 sky130_fd_sc_hd__or2b_2 _23641_ (.A(_13162_),
    .B_N(_13161_),
    .X(_13418_));
 sky130_fd_sc_hd__and4_2 _23642_ (.A(iX[13]),
    .B(iX[14]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_13419_));
 sky130_fd_sc_hd__a22oi_2 _23643_ (.A1(iX[14]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[13]),
    .Y(_13421_));
 sky130_fd_sc_hd__nor2_2 _23644_ (.A(_13419_),
    .B(_13421_),
    .Y(_13422_));
 sky130_fd_sc_hd__nand2_2 _23645_ (.A(iX[12]),
    .B(iY[29]),
    .Y(_13423_));
 sky130_fd_sc_hd__xnor2_2 _23646_ (.A(_13422_),
    .B(_13423_),
    .Y(_13424_));
 sky130_fd_sc_hd__o21ba_2 _23647_ (.A1(_13157_),
    .A2(_13160_),
    .B1_N(_13156_),
    .X(_13425_));
 sky130_fd_sc_hd__xnor2_2 _23648_ (.A(_13424_),
    .B(_13425_),
    .Y(_13426_));
 sky130_fd_sc_hd__nand3_2 _23649_ (.A(iX[11]),
    .B(iY[30]),
    .C(_13426_),
    .Y(_13427_));
 sky130_fd_sc_hd__a21o_2 _23650_ (.A1(iX[11]),
    .A2(iY[30]),
    .B1(_13426_),
    .X(_13428_));
 sky130_fd_sc_hd__nand2_2 _23651_ (.A(_13427_),
    .B(_13428_),
    .Y(_13429_));
 sky130_fd_sc_hd__a21oi_2 _23652_ (.A1(_13418_),
    .A2(_13164_),
    .B1(_13429_),
    .Y(_13430_));
 sky130_fd_sc_hd__and3_2 _23653_ (.A(_13418_),
    .B(_13164_),
    .C(_13429_),
    .X(_13432_));
 sky130_fd_sc_hd__nor2_2 _23654_ (.A(_13430_),
    .B(_13432_),
    .Y(_13433_));
 sky130_fd_sc_hd__a21oi_2 _23655_ (.A1(iX[10]),
    .A2(iY[31]),
    .B1(_13433_),
    .Y(_13434_));
 sky130_fd_sc_hd__and3_2 _23656_ (.A(iX[10]),
    .B(iY[31]),
    .C(_13433_),
    .X(_13435_));
 sky130_fd_sc_hd__nor2_2 _23657_ (.A(_13434_),
    .B(_13435_),
    .Y(_13436_));
 sky130_fd_sc_hd__or2b_2 _23658_ (.A(_13179_),
    .B_N(_13185_),
    .X(_13437_));
 sky130_fd_sc_hd__or2b_2 _23659_ (.A(_13178_),
    .B_N(_13186_),
    .X(_13438_));
 sky130_fd_sc_hd__and2b_2 _23660_ (.A_N(_13121_),
    .B(_13120_),
    .X(_13439_));
 sky130_fd_sc_hd__o21ba_2 _23661_ (.A1(_13182_),
    .A2(_13184_),
    .B1_N(_13181_),
    .X(_13440_));
 sky130_fd_sc_hd__o21ba_2 _23662_ (.A1(_13111_),
    .A2(_13113_),
    .B1_N(_13110_),
    .X(_13441_));
 sky130_fd_sc_hd__and4_2 _23663_ (.A(iX[16]),
    .B(iX[17]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_13443_));
 sky130_fd_sc_hd__a22oi_2 _23664_ (.A1(iX[17]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[16]),
    .Y(_13444_));
 sky130_fd_sc_hd__nor2_2 _23665_ (.A(_13443_),
    .B(_13444_),
    .Y(_13445_));
 sky130_fd_sc_hd__nand2_2 _23666_ (.A(iX[15]),
    .B(iY[26]),
    .Y(_13446_));
 sky130_fd_sc_hd__xnor2_2 _23667_ (.A(_13445_),
    .B(_13446_),
    .Y(_13447_));
 sky130_fd_sc_hd__xnor2_2 _23668_ (.A(_13441_),
    .B(_13447_),
    .Y(_13448_));
 sky130_fd_sc_hd__xnor2_2 _23669_ (.A(_13440_),
    .B(_13448_),
    .Y(_13449_));
 sky130_fd_sc_hd__o21a_2 _23670_ (.A1(_13439_),
    .A2(_13123_),
    .B1(_13449_),
    .X(_13450_));
 sky130_fd_sc_hd__nor3_2 _23671_ (.A(_13439_),
    .B(_13123_),
    .C(_13449_),
    .Y(_13451_));
 sky130_fd_sc_hd__a211oi_2 _23672_ (.A1(_13437_),
    .A2(_13438_),
    .B1(_13450_),
    .C1(_13451_),
    .Y(_13452_));
 sky130_fd_sc_hd__o211a_2 _23673_ (.A1(_13450_),
    .A2(_13451_),
    .B1(_13437_),
    .C1(_13438_),
    .X(_13454_));
 sky130_fd_sc_hd__nor2_2 _23674_ (.A(_13188_),
    .B(_13190_),
    .Y(_13455_));
 sky130_fd_sc_hd__or3_2 _23675_ (.A(_13452_),
    .B(_13454_),
    .C(_13455_),
    .X(_13456_));
 sky130_fd_sc_hd__o21ai_2 _23676_ (.A1(_13452_),
    .A2(_13454_),
    .B1(_13455_),
    .Y(_13457_));
 sky130_fd_sc_hd__and3_2 _23677_ (.A(_13436_),
    .B(_13456_),
    .C(_13457_),
    .X(_13458_));
 sky130_fd_sc_hd__a21oi_2 _23678_ (.A1(_13456_),
    .A2(_13457_),
    .B1(_13436_),
    .Y(_13459_));
 sky130_fd_sc_hd__or3_2 _23679_ (.A(_13417_),
    .B(_13458_),
    .C(_13459_),
    .X(_13460_));
 sky130_fd_sc_hd__o21ai_2 _23680_ (.A1(_13458_),
    .A2(_13459_),
    .B1(_13417_),
    .Y(_13461_));
 sky130_fd_sc_hd__nand2_2 _23681_ (.A(_13460_),
    .B(_13461_),
    .Y(_13462_));
 sky130_fd_sc_hd__a21o_2 _23682_ (.A1(_13194_),
    .A2(_13415_),
    .B1(_13462_),
    .X(_13463_));
 sky130_fd_sc_hd__nand3_2 _23683_ (.A(_13194_),
    .B(_13415_),
    .C(_13462_),
    .Y(_13465_));
 sky130_fd_sc_hd__nand4_2 _23684_ (.A(_13413_),
    .B(_13414_),
    .C(_13463_),
    .D(_13465_),
    .Y(_13466_));
 sky130_fd_sc_hd__a22o_2 _23685_ (.A1(_13413_),
    .A2(_13414_),
    .B1(_13463_),
    .B2(_13465_),
    .X(_13467_));
 sky130_fd_sc_hd__nand2_2 _23686_ (.A(_13151_),
    .B(_13204_),
    .Y(_13468_));
 sky130_fd_sc_hd__and3_2 _23687_ (.A(_13466_),
    .B(_13467_),
    .C(_13468_),
    .X(_13469_));
 sky130_fd_sc_hd__a21oi_2 _23688_ (.A1(_13466_),
    .A2(_13467_),
    .B1(_13468_),
    .Y(_13470_));
 sky130_fd_sc_hd__a211oi_2 _23689_ (.A1(_13198_),
    .A2(_13201_),
    .B1(_13469_),
    .C1(_13470_),
    .Y(_13471_));
 sky130_fd_sc_hd__o211a_2 _23690_ (.A1(_13469_),
    .A2(_13470_),
    .B1(_13198_),
    .C1(_13201_),
    .X(_13472_));
 sky130_fd_sc_hd__nor2_2 _23691_ (.A(_13471_),
    .B(_13472_),
    .Y(_13473_));
 sky130_fd_sc_hd__o21a_2 _23692_ (.A1(_13206_),
    .A2(_13351_),
    .B1(_13473_),
    .X(_13474_));
 sky130_fd_sc_hd__nor3_2 _23693_ (.A(_13206_),
    .B(_13351_),
    .C(_13473_),
    .Y(_13476_));
 sky130_fd_sc_hd__inv_2 _23694_ (.A(_13166_),
    .Y(_13477_));
 sky130_fd_sc_hd__a21oi_2 _23695_ (.A1(_13477_),
    .A2(_13168_),
    .B1(_13173_),
    .Y(_13478_));
 sky130_fd_sc_hd__nor3_2 _23696_ (.A(_13474_),
    .B(_13476_),
    .C(_13478_),
    .Y(_13479_));
 sky130_fd_sc_hd__o21a_2 _23697_ (.A1(_13474_),
    .A2(_13476_),
    .B1(_13478_),
    .X(_13480_));
 sky130_fd_sc_hd__or2_2 _23698_ (.A(_13479_),
    .B(_13480_),
    .X(_13481_));
 sky130_fd_sc_hd__a21oi_2 _23699_ (.A1(_13214_),
    .A2(_13215_),
    .B1(_13211_),
    .Y(_13482_));
 sky130_fd_sc_hd__xnor2_2 _23700_ (.A(_13481_),
    .B(_13482_),
    .Y(_13483_));
 sky130_fd_sc_hd__nor2_2 _23701_ (.A(_13218_),
    .B(_13483_),
    .Y(_13484_));
 sky130_fd_sc_hd__a311o_2 _23702_ (.A1(_12204_),
    .A2(_12209_),
    .A3(_13225_),
    .B1(_13227_),
    .C1(_13220_),
    .X(_13485_));
 sky130_fd_sc_hd__nor2_2 _23703_ (.A(_13485_),
    .B(_13483_),
    .Y(_13487_));
 sky130_fd_sc_hd__and3_2 _23704_ (.A(_13218_),
    .B(_13485_),
    .C(_13483_),
    .X(_13488_));
 sky130_fd_sc_hd__or3_2 _23705_ (.A(_13484_),
    .B(_13487_),
    .C(_13488_),
    .X(_13489_));
 sky130_fd_sc_hd__a211o_2 _23706_ (.A1(_12858_),
    .A2(_12860_),
    .B1(_13286_),
    .C1(_13287_),
    .X(_13490_));
 sky130_fd_sc_hd__and2_2 _23707_ (.A(iX[9]),
    .B(iX[41]),
    .X(_13491_));
 sky130_fd_sc_hd__nor2_2 _23708_ (.A(iX[9]),
    .B(iX[41]),
    .Y(_13492_));
 sky130_fd_sc_hd__or2_2 _23709_ (.A(_13491_),
    .B(_13492_),
    .X(_13493_));
 sky130_fd_sc_hd__buf_1 _23710_ (.A(_13493_),
    .X(_13494_));
 sky130_fd_sc_hd__a21oi_4 _23711_ (.A1(_13237_),
    .A2(_13240_),
    .B1(_13238_),
    .Y(_13495_));
 sky130_fd_sc_hd__xor2_2 _23712_ (.A(_13494_),
    .B(_13495_),
    .X(_13496_));
 sky130_fd_sc_hd__and3_2 _23713_ (.A(_11378_),
    .B(_13242_),
    .C(_13496_),
    .X(_13498_));
 sky130_fd_sc_hd__a21o_2 _23714_ (.A1(_11379_),
    .A2(_13496_),
    .B1(_13242_),
    .X(_13499_));
 sky130_fd_sc_hd__or4b_4 _23715_ (.A(_11791_),
    .B(_12808_),
    .C(_13498_),
    .D_N(_13499_),
    .X(_13500_));
 sky130_fd_sc_hd__buf_1 _23716_ (.A(_12811_),
    .X(_13501_));
 sky130_fd_sc_hd__xnor2_2 _23717_ (.A(_13494_),
    .B(_13495_),
    .Y(_13502_));
 sky130_fd_sc_hd__or3b_2 _23718_ (.A(_11565_),
    .B(_13502_),
    .C_N(_13242_),
    .X(_13503_));
 sky130_fd_sc_hd__a22o_2 _23719_ (.A1(_12450_),
    .A2(_13501_),
    .B1(_13503_),
    .B2(_13499_),
    .X(_13504_));
 sky130_fd_sc_hd__a31o_2 _23720_ (.A1(_12450_),
    .A2(_12816_),
    .A3(_13245_),
    .B1(_13243_),
    .X(_13505_));
 sky130_fd_sc_hd__nand3_2 _23721_ (.A(_13500_),
    .B(_13504_),
    .C(_13505_),
    .Y(_13506_));
 sky130_fd_sc_hd__a21o_2 _23722_ (.A1(_13500_),
    .A2(_13504_),
    .B1(_13505_),
    .X(_13507_));
 sky130_fd_sc_hd__and3_2 _23723_ (.A(_12241_),
    .B(_12810_),
    .C(_13253_),
    .X(_13509_));
 sky130_fd_sc_hd__o22a_2 _23724_ (.A1(_12247_),
    .A2(_12457_),
    .B1(_13231_),
    .B2(_12244_),
    .X(_13510_));
 sky130_fd_sc_hd__nor2_2 _23725_ (.A(_13509_),
    .B(_13510_),
    .Y(_13511_));
 sky130_fd_sc_hd__nand2_2 _23726_ (.A(_12225_),
    .B(_12477_),
    .Y(_13512_));
 sky130_fd_sc_hd__xnor2_2 _23727_ (.A(_13511_),
    .B(_13512_),
    .Y(_13513_));
 sky130_fd_sc_hd__nand3_2 _23728_ (.A(_13506_),
    .B(_13507_),
    .C(_13513_),
    .Y(_13514_));
 sky130_fd_sc_hd__a21o_2 _23729_ (.A1(_13506_),
    .A2(_13507_),
    .B1(_13513_),
    .X(_13515_));
 sky130_fd_sc_hd__a21bo_2 _23730_ (.A1(_13252_),
    .A2(_13256_),
    .B1_N(_13251_),
    .X(_13516_));
 sky130_fd_sc_hd__and3_2 _23731_ (.A(_13514_),
    .B(_13515_),
    .C(_13516_),
    .X(_13517_));
 sky130_fd_sc_hd__a21oi_2 _23732_ (.A1(_13514_),
    .A2(_13515_),
    .B1(_13516_),
    .Y(_13518_));
 sky130_fd_sc_hd__nand2_2 _23733_ (.A(_13265_),
    .B(_13275_),
    .Y(_13520_));
 sky130_fd_sc_hd__and3_2 _23734_ (.A(_11829_),
    .B(_12477_),
    .C(_13254_),
    .X(_13521_));
 sky130_fd_sc_hd__a31o_2 _23735_ (.A1(_12225_),
    .A2(_12242_),
    .A3(_13253_),
    .B1(_13521_),
    .X(_13522_));
 sky130_fd_sc_hd__and3_2 _23736_ (.A(_11829_),
    .B(_12845_),
    .C(_13264_),
    .X(_13523_));
 sky130_fd_sc_hd__o22a_2 _23737_ (.A1(_11827_),
    .A2(_12772_),
    .B1(_12849_),
    .B2(_12468_),
    .X(_13524_));
 sky130_fd_sc_hd__or4_2 _23738_ (.A(_11569_),
    .B(_13273_),
    .C(_13523_),
    .D(_13524_),
    .X(_13525_));
 sky130_fd_sc_hd__a2bb2o_2 _23739_ (.A1_N(_13523_),
    .A2_N(_13524_),
    .B1(_11581_),
    .B2(_13274_),
    .X(_13526_));
 sky130_fd_sc_hd__nand3_2 _23740_ (.A(_13522_),
    .B(_13525_),
    .C(_13526_),
    .Y(_13527_));
 sky130_fd_sc_hd__a21o_2 _23741_ (.A1(_13525_),
    .A2(_13526_),
    .B1(_13522_),
    .X(_13528_));
 sky130_fd_sc_hd__and3_2 _23742_ (.A(_13520_),
    .B(_13527_),
    .C(_13528_),
    .X(_13529_));
 sky130_fd_sc_hd__a21oi_2 _23743_ (.A1(_13527_),
    .A2(_13528_),
    .B1(_13520_),
    .Y(_13531_));
 sky130_fd_sc_hd__nor4_2 _23744_ (.A(_13517_),
    .B(_13518_),
    .C(_13529_),
    .D(_13531_),
    .Y(_13532_));
 sky130_fd_sc_hd__o22a_2 _23745_ (.A1(_13517_),
    .A2(_13518_),
    .B1(_13529_),
    .B2(_13531_),
    .X(_13533_));
 sky130_fd_sc_hd__a211oi_2 _23746_ (.A1(_13261_),
    .A2(_13282_),
    .B1(_13532_),
    .C1(_13533_),
    .Y(_13534_));
 sky130_fd_sc_hd__o211a_2 _23747_ (.A1(_13532_),
    .A2(_13533_),
    .B1(_13261_),
    .C1(_13282_),
    .X(_13535_));
 sky130_fd_sc_hd__or2_4 _23748_ (.A(iY[9]),
    .B(iY[41]),
    .X(_13536_));
 sky130_fd_sc_hd__nand2_2 _23749_ (.A(iY[9]),
    .B(iY[41]),
    .Y(_13537_));
 sky130_fd_sc_hd__and2_2 _23750_ (.A(_13536_),
    .B(_13537_),
    .X(_13538_));
 sky130_fd_sc_hd__o211a_2 _23751_ (.A1(_12771_),
    .A2(_13269_),
    .B1(_13271_),
    .C1(_13267_),
    .X(_13539_));
 sky130_fd_sc_hd__a21o_2 _23752_ (.A1(iY[8]),
    .A2(iY[40]),
    .B1(_13539_),
    .X(_13540_));
 sky130_fd_sc_hd__xor2_2 _23753_ (.A(_13538_),
    .B(_13540_),
    .X(_13542_));
 sky130_fd_sc_hd__buf_1 _23754_ (.A(_13542_),
    .X(_13543_));
 sky130_fd_sc_hd__buf_1 _23755_ (.A(_13543_),
    .X(_13544_));
 sky130_fd_sc_hd__nand2_2 _23756_ (.A(_11374_),
    .B(_13544_),
    .Y(_13545_));
 sky130_fd_sc_hd__a21oi_2 _23757_ (.A1(_13277_),
    .A2(_13281_),
    .B1(_13545_),
    .Y(_13546_));
 sky130_fd_sc_hd__and3_2 _23758_ (.A(_13277_),
    .B(_13281_),
    .C(_13545_),
    .X(_13547_));
 sky130_fd_sc_hd__or2_2 _23759_ (.A(_13546_),
    .B(_13547_),
    .X(_13548_));
 sky130_fd_sc_hd__or3_2 _23760_ (.A(_13534_),
    .B(_13535_),
    .C(_13548_),
    .X(_13549_));
 sky130_fd_sc_hd__o21ai_2 _23761_ (.A1(_13534_),
    .A2(_13535_),
    .B1(_13548_),
    .Y(_13550_));
 sky130_fd_sc_hd__o211a_2 _23762_ (.A1(_13284_),
    .A2(_13286_),
    .B1(_13549_),
    .C1(_13550_),
    .X(_13551_));
 sky130_fd_sc_hd__a211oi_2 _23763_ (.A1(_13549_),
    .A2(_13550_),
    .B1(_13284_),
    .C1(_13286_),
    .Y(_13553_));
 sky130_fd_sc_hd__nor3_2 _23764_ (.A(_13490_),
    .B(_13551_),
    .C(_13553_),
    .Y(_13554_));
 sky130_fd_sc_hd__o21a_2 _23765_ (.A1(_13551_),
    .A2(_13553_),
    .B1(_13490_),
    .X(_13555_));
 sky130_fd_sc_hd__and4bb_2 _23766_ (.A_N(_13554_),
    .B_N(_13555_),
    .C(_12863_),
    .D(_13291_),
    .X(_13556_));
 sky130_fd_sc_hd__o2bb2a_2 _23767_ (.A1_N(_12863_),
    .A2_N(_13291_),
    .B1(_13554_),
    .B2(_13555_),
    .X(_13557_));
 sky130_fd_sc_hd__nor2_2 _23768_ (.A(_12784_),
    .B(_13294_),
    .Y(_13558_));
 sky130_fd_sc_hd__or4bb_4 _23769_ (.A(_13556_),
    .B(_13557_),
    .C_N(_13291_),
    .D_N(_13558_),
    .X(_13559_));
 sky130_fd_sc_hd__a2bb2o_2 _23770_ (.A1_N(_13556_),
    .A2_N(_13557_),
    .B1(_13291_),
    .B2(_13558_),
    .X(_13560_));
 sky130_fd_sc_hd__and2_2 _23771_ (.A(_13293_),
    .B(_13295_),
    .X(_13561_));
 sky130_fd_sc_hd__a21oi_2 _23772_ (.A1(_13559_),
    .A2(_13560_),
    .B1(_13561_),
    .Y(_13562_));
 sky130_fd_sc_hd__and3_2 _23773_ (.A(_13561_),
    .B(_13559_),
    .C(_13560_),
    .X(_13564_));
 sky130_fd_sc_hd__or2_2 _23774_ (.A(_12902_),
    .B(_13335_),
    .X(_13565_));
 sky130_fd_sc_hd__nand2_2 _23775_ (.A(_13333_),
    .B(_13334_),
    .Y(_13566_));
 sky130_fd_sc_hd__and4_2 _23776_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[38]),
    .D(iX[39]),
    .X(_13567_));
 sky130_fd_sc_hd__a22oi_2 _23777_ (.A1(iY[35]),
    .A2(iX[38]),
    .B1(iX[39]),
    .B2(iY[34]),
    .Y(_13568_));
 sky130_fd_sc_hd__nand2_2 _23778_ (.A(iY[33]),
    .B(iX[40]),
    .Y(_13569_));
 sky130_fd_sc_hd__or3_2 _23779_ (.A(_13567_),
    .B(_13568_),
    .C(_13569_),
    .X(_13570_));
 sky130_fd_sc_hd__o21ai_2 _23780_ (.A1(_13567_),
    .A2(_13568_),
    .B1(_13569_),
    .Y(_13571_));
 sky130_fd_sc_hd__o21bai_2 _23781_ (.A1(_13299_),
    .A2(_13300_),
    .B1_N(_13298_),
    .Y(_13572_));
 sky130_fd_sc_hd__nand3_2 _23782_ (.A(_13570_),
    .B(_13571_),
    .C(_13572_),
    .Y(_13573_));
 sky130_fd_sc_hd__a21o_2 _23783_ (.A1(_13570_),
    .A2(_13571_),
    .B1(_13572_),
    .X(_13575_));
 sky130_fd_sc_hd__and4_2 _23784_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[37]),
    .D(iX[41]),
    .X(_13576_));
 sky130_fd_sc_hd__a22oi_2 _23785_ (.A1(iY[36]),
    .A2(iX[37]),
    .B1(iX[41]),
    .B2(iY[32]),
    .Y(_13577_));
 sky130_fd_sc_hd__nor2_2 _23786_ (.A(_13576_),
    .B(_13577_),
    .Y(_13578_));
 sky130_fd_sc_hd__nand2_2 _23787_ (.A(iX[36]),
    .B(iY[37]),
    .Y(_13579_));
 sky130_fd_sc_hd__xnor2_2 _23788_ (.A(_13578_),
    .B(_13579_),
    .Y(_13580_));
 sky130_fd_sc_hd__nand3_2 _23789_ (.A(_13573_),
    .B(_13575_),
    .C(_13580_),
    .Y(_13581_));
 sky130_fd_sc_hd__a21o_2 _23790_ (.A1(_13573_),
    .A2(_13575_),
    .B1(_13580_),
    .X(_13582_));
 sky130_fd_sc_hd__a21bo_2 _23791_ (.A1(_13306_),
    .A2(_13311_),
    .B1_N(_13305_),
    .X(_13583_));
 sky130_fd_sc_hd__nand3_2 _23792_ (.A(_13581_),
    .B(_13582_),
    .C(_13583_),
    .Y(_13584_));
 sky130_fd_sc_hd__a21o_2 _23793_ (.A1(_13581_),
    .A2(_13582_),
    .B1(_13583_),
    .X(_13586_));
 sky130_fd_sc_hd__o21ba_2 _23794_ (.A1(_13320_),
    .A2(_13322_),
    .B1_N(_13319_),
    .X(_13587_));
 sky130_fd_sc_hd__o21ba_2 _23795_ (.A1(_13308_),
    .A2(_13310_),
    .B1_N(_13307_),
    .X(_13588_));
 sky130_fd_sc_hd__and4_2 _23796_ (.A(iX[34]),
    .B(iX[35]),
    .C(iY[38]),
    .D(iY[39]),
    .X(_13589_));
 sky130_fd_sc_hd__a22oi_2 _23797_ (.A1(iX[35]),
    .A2(iY[38]),
    .B1(iY[39]),
    .B2(iX[34]),
    .Y(_13590_));
 sky130_fd_sc_hd__nor2_2 _23798_ (.A(_13589_),
    .B(_13590_),
    .Y(_13591_));
 sky130_fd_sc_hd__nand2_2 _23799_ (.A(iX[33]),
    .B(iY[40]),
    .Y(_13592_));
 sky130_fd_sc_hd__xnor2_2 _23800_ (.A(_13591_),
    .B(_13592_),
    .Y(_13593_));
 sky130_fd_sc_hd__xnor2_2 _23801_ (.A(_13588_),
    .B(_13593_),
    .Y(_13594_));
 sky130_fd_sc_hd__xnor2_2 _23802_ (.A(_13587_),
    .B(_13594_),
    .Y(_13595_));
 sky130_fd_sc_hd__nand3_2 _23803_ (.A(_13584_),
    .B(_13586_),
    .C(_13595_),
    .Y(_13597_));
 sky130_fd_sc_hd__a21o_2 _23804_ (.A1(_13584_),
    .A2(_13586_),
    .B1(_13595_),
    .X(_13598_));
 sky130_fd_sc_hd__o211a_2 _23805_ (.A1(_13316_),
    .A2(_13327_),
    .B1(_13597_),
    .C1(_13598_),
    .X(_13599_));
 sky130_fd_sc_hd__a211o_2 _23806_ (.A1(_13597_),
    .A2(_13598_),
    .B1(_13316_),
    .C1(_13327_),
    .X(_13600_));
 sky130_fd_sc_hd__or2b_2 _23807_ (.A(_13599_),
    .B_N(_13600_),
    .X(_13601_));
 sky130_fd_sc_hd__and2_2 _23808_ (.A(_13318_),
    .B(_13324_),
    .X(_13602_));
 sky130_fd_sc_hd__and2_2 _23809_ (.A(_12888_),
    .B(_13325_),
    .X(_13603_));
 sky130_fd_sc_hd__o211a_2 _23810_ (.A1(_13602_),
    .A2(_13603_),
    .B1(iX[32]),
    .C1(iY[41]),
    .X(_13604_));
 sky130_fd_sc_hd__a211oi_2 _23811_ (.A1(iX[32]),
    .A2(iY[41]),
    .B1(_13602_),
    .C1(_13603_),
    .Y(_13605_));
 sky130_fd_sc_hd__nor2_2 _23812_ (.A(_13604_),
    .B(_13605_),
    .Y(_13606_));
 sky130_fd_sc_hd__xnor2_2 _23813_ (.A(_13601_),
    .B(_13606_),
    .Y(_13608_));
 sky130_fd_sc_hd__or2_2 _23814_ (.A(_13329_),
    .B(_13332_),
    .X(_13609_));
 sky130_fd_sc_hd__xnor2_2 _23815_ (.A(_13608_),
    .B(_13609_),
    .Y(_13610_));
 sky130_fd_sc_hd__xor2_2 _23816_ (.A(_13566_),
    .B(_13610_),
    .X(_13611_));
 sky130_fd_sc_hd__xnor2_2 _23817_ (.A(_13565_),
    .B(_13611_),
    .Y(_13612_));
 sky130_fd_sc_hd__or3_2 _23818_ (.A(_12905_),
    .B(_12904_),
    .C(_13335_),
    .X(_13613_));
 sky130_fd_sc_hd__o31a_2 _23819_ (.A1(_12733_),
    .A2(_12904_),
    .A3(_13337_),
    .B1(_13613_),
    .X(_13614_));
 sky130_fd_sc_hd__xnor2_2 _23820_ (.A(_13612_),
    .B(_13614_),
    .Y(_13615_));
 sky130_fd_sc_hd__xor2_2 _23821_ (.A(_13339_),
    .B(_13615_),
    .X(_13616_));
 sky130_fd_sc_hd__nor3_2 _23822_ (.A(_13562_),
    .B(_13564_),
    .C(_13616_),
    .Y(_13617_));
 sky130_fd_sc_hd__o21a_2 _23823_ (.A1(_13562_),
    .A2(_13564_),
    .B1(_13616_),
    .X(_13619_));
 sky130_fd_sc_hd__or3_2 _23824_ (.A(oO[9]),
    .B(_13617_),
    .C(_13619_),
    .X(_13620_));
 sky130_fd_sc_hd__o21ai_2 _23825_ (.A1(_13617_),
    .A2(_13619_),
    .B1(oO[9]),
    .Y(_13621_));
 sky130_fd_sc_hd__or2_2 _23826_ (.A(_13296_),
    .B(_13341_),
    .X(_13622_));
 sky130_fd_sc_hd__o21ai_2 _23827_ (.A1(oO[8]),
    .A2(_13342_),
    .B1(_13622_),
    .Y(_13623_));
 sky130_fd_sc_hd__and3_2 _23828_ (.A(_13620_),
    .B(_13621_),
    .C(_13623_),
    .X(_13624_));
 sky130_fd_sc_hd__a21oi_2 _23829_ (.A1(_13620_),
    .A2(_13621_),
    .B1(_13623_),
    .Y(_13625_));
 sky130_fd_sc_hd__or2_2 _23830_ (.A(_13624_),
    .B(_13625_),
    .X(_13626_));
 sky130_fd_sc_hd__or2b_2 _23831_ (.A(_13346_),
    .B_N(_13348_),
    .X(_13627_));
 sky130_fd_sc_hd__o21a_2 _23832_ (.A1(_13343_),
    .A2(_13345_),
    .B1(_13627_),
    .X(_13628_));
 sky130_fd_sc_hd__xor2_2 _23833_ (.A(_13626_),
    .B(_13628_),
    .X(_13630_));
 sky130_fd_sc_hd__and2b_2 _23834_ (.A_N(_13489_),
    .B(_13630_),
    .X(_13631_));
 sky130_fd_sc_hd__and2b_2 _23835_ (.A_N(_13630_),
    .B(_13489_),
    .X(_13632_));
 sky130_fd_sc_hd__or2_2 _23836_ (.A(_13631_),
    .B(_13632_),
    .X(_13633_));
 sky130_fd_sc_hd__and2b_2 _23837_ (.A_N(_13229_),
    .B(_13349_),
    .X(_13634_));
 sky130_fd_sc_hd__a21o_2 _23838_ (.A1(_13073_),
    .A2(_13350_),
    .B1(_13634_),
    .X(_13635_));
 sky130_fd_sc_hd__xnor2_2 _23839_ (.A(_13633_),
    .B(_13635_),
    .Y(oO[41]));
 sky130_fd_sc_hd__or3b_2 _23840_ (.A(_13631_),
    .B(_13632_),
    .C_N(_13350_),
    .X(_13636_));
 sky130_fd_sc_hd__a21oi_2 _23841_ (.A1(_13071_),
    .A2(_13072_),
    .B1(_13636_),
    .Y(_13637_));
 sky130_fd_sc_hd__o21ba_2 _23842_ (.A1(_13634_),
    .A2(_13631_),
    .B1_N(_13632_),
    .X(_13638_));
 sky130_fd_sc_hd__or2_2 _23843_ (.A(_13637_),
    .B(_13638_),
    .X(_13640_));
 sky130_fd_sc_hd__or2b_2 _23844_ (.A(_13356_),
    .B_N(_13357_),
    .X(_13641_));
 sky130_fd_sc_hd__and3b_2 _23845_ (.A_N(_12932_),
    .B(iX[31]),
    .C(iY[11]),
    .X(_13642_));
 sky130_fd_sc_hd__and2_2 _23846_ (.A(iY[13]),
    .B(iX[30]),
    .X(_13643_));
 sky130_fd_sc_hd__and3_2 _23847_ (.A(iY[12]),
    .B(iX[29]),
    .C(_13643_),
    .X(_13644_));
 sky130_fd_sc_hd__a22oi_2 _23848_ (.A1(iY[13]),
    .A2(iX[29]),
    .B1(iX[30]),
    .B2(iY[12]),
    .Y(_13645_));
 sky130_fd_sc_hd__and4bb_2 _23849_ (.A_N(_13644_),
    .B_N(_13645_),
    .C(iY[14]),
    .D(iX[28]),
    .X(_13646_));
 sky130_fd_sc_hd__o2bb2a_2 _23850_ (.A1_N(iY[14]),
    .A2_N(iX[28]),
    .B1(_13644_),
    .B2(_13645_),
    .X(_13647_));
 sky130_fd_sc_hd__nor2_2 _23851_ (.A(_13646_),
    .B(_13647_),
    .Y(_13648_));
 sky130_fd_sc_hd__xnor2_2 _23852_ (.A(_13642_),
    .B(_13648_),
    .Y(_13649_));
 sky130_fd_sc_hd__a21oi_2 _23853_ (.A1(_13641_),
    .A2(_13364_),
    .B1(_13649_),
    .Y(_13651_));
 sky130_fd_sc_hd__and3_2 _23854_ (.A(_13641_),
    .B(_13364_),
    .C(_13649_),
    .X(_13652_));
 sky130_fd_sc_hd__or2_2 _23855_ (.A(_13651_),
    .B(_13652_),
    .X(_13653_));
 sky130_fd_sc_hd__a21o_2 _23856_ (.A1(_13390_),
    .A2(_13135_),
    .B1(_13401_),
    .X(_13654_));
 sky130_fd_sc_hd__and4_2 _23857_ (.A(iX[20]),
    .B(iX[21]),
    .C(iY[21]),
    .D(iY[22]),
    .X(_13655_));
 sky130_fd_sc_hd__a22oi_2 _23858_ (.A1(iX[21]),
    .A2(iY[21]),
    .B1(iY[22]),
    .B2(iX[20]),
    .Y(_13656_));
 sky130_fd_sc_hd__nor2_2 _23859_ (.A(_13655_),
    .B(_13656_),
    .Y(_13657_));
 sky130_fd_sc_hd__nand2_2 _23860_ (.A(iX[19]),
    .B(iY[23]),
    .Y(_13658_));
 sky130_fd_sc_hd__xnor2_2 _23861_ (.A(_13657_),
    .B(_13658_),
    .Y(_13659_));
 sky130_fd_sc_hd__and4_2 _23862_ (.A(iY[18]),
    .B(iY[19]),
    .C(iX[23]),
    .D(iX[24]),
    .X(_13660_));
 sky130_fd_sc_hd__a22oi_2 _23863_ (.A1(iY[19]),
    .A2(iX[23]),
    .B1(iX[24]),
    .B2(iY[18]),
    .Y(_13662_));
 sky130_fd_sc_hd__nor2_2 _23864_ (.A(_13660_),
    .B(_13662_),
    .Y(_13663_));
 sky130_fd_sc_hd__nand2_2 _23865_ (.A(iY[20]),
    .B(iX[22]),
    .Y(_13664_));
 sky130_fd_sc_hd__xnor2_2 _23866_ (.A(_13663_),
    .B(_13664_),
    .Y(_13665_));
 sky130_fd_sc_hd__o21ba_2 _23867_ (.A1(_13380_),
    .A2(_13382_),
    .B1_N(_13379_),
    .X(_13666_));
 sky130_fd_sc_hd__xnor2_2 _23868_ (.A(_13665_),
    .B(_13666_),
    .Y(_13667_));
 sky130_fd_sc_hd__and2_2 _23869_ (.A(_13659_),
    .B(_13667_),
    .X(_13668_));
 sky130_fd_sc_hd__nor2_2 _23870_ (.A(_13659_),
    .B(_13667_),
    .Y(_13669_));
 sky130_fd_sc_hd__or2_2 _23871_ (.A(_13668_),
    .B(_13669_),
    .X(_13670_));
 sky130_fd_sc_hd__nand2_2 _23872_ (.A(_13391_),
    .B(_13400_),
    .Y(_13671_));
 sky130_fd_sc_hd__o21ba_2 _23873_ (.A1(_13360_),
    .A2(_13362_),
    .B1_N(_13359_),
    .X(_13673_));
 sky130_fd_sc_hd__and4_2 _23874_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[26]),
    .D(iX[27]),
    .X(_13674_));
 sky130_fd_sc_hd__a22oi_2 _23875_ (.A1(iY[16]),
    .A2(iX[26]),
    .B1(iX[27]),
    .B2(iY[15]),
    .Y(_13675_));
 sky130_fd_sc_hd__nor2_2 _23876_ (.A(_13674_),
    .B(_13675_),
    .Y(_13676_));
 sky130_fd_sc_hd__nand2_2 _23877_ (.A(iY[17]),
    .B(iX[25]),
    .Y(_13677_));
 sky130_fd_sc_hd__xnor2_2 _23878_ (.A(_13676_),
    .B(_13677_),
    .Y(_13678_));
 sky130_fd_sc_hd__xnor2_2 _23879_ (.A(_13673_),
    .B(_13678_),
    .Y(_13679_));
 sky130_fd_sc_hd__o21ai_2 _23880_ (.A1(_13392_),
    .A2(_13394_),
    .B1(_13679_),
    .Y(_13680_));
 sky130_fd_sc_hd__or3_2 _23881_ (.A(_13392_),
    .B(_13394_),
    .C(_13679_),
    .X(_13681_));
 sky130_fd_sc_hd__nand2_2 _23882_ (.A(_13680_),
    .B(_13681_),
    .Y(_13682_));
 sky130_fd_sc_hd__a21oi_2 _23883_ (.A1(_13397_),
    .A2(_13671_),
    .B1(_13682_),
    .Y(_13684_));
 sky130_fd_sc_hd__and3_2 _23884_ (.A(_13397_),
    .B(_13671_),
    .C(_13682_),
    .X(_13685_));
 sky130_fd_sc_hd__or3_2 _23885_ (.A(_13670_),
    .B(_13684_),
    .C(_13685_),
    .X(_13686_));
 sky130_fd_sc_hd__o21ai_2 _23886_ (.A1(_13684_),
    .A2(_13685_),
    .B1(_13670_),
    .Y(_13687_));
 sky130_fd_sc_hd__and3_2 _23887_ (.A(_13368_),
    .B(_13686_),
    .C(_13687_),
    .X(_13688_));
 sky130_fd_sc_hd__a21oi_2 _23888_ (.A1(_13686_),
    .A2(_13687_),
    .B1(_13368_),
    .Y(_13689_));
 sky130_fd_sc_hd__a211oi_2 _23889_ (.A1(_13654_),
    .A2(_13404_),
    .B1(_13688_),
    .C1(_13689_),
    .Y(_13690_));
 sky130_fd_sc_hd__o211a_2 _23890_ (.A1(_13688_),
    .A2(_13689_),
    .B1(_13654_),
    .C1(_13404_),
    .X(_13691_));
 sky130_fd_sc_hd__or3_2 _23891_ (.A(_13653_),
    .B(_13690_),
    .C(_13691_),
    .X(_13692_));
 sky130_fd_sc_hd__inv_2 _23892_ (.A(_13692_),
    .Y(_13693_));
 sky130_fd_sc_hd__o21a_2 _23893_ (.A1(_13690_),
    .A2(_13691_),
    .B1(_13653_),
    .X(_13695_));
 sky130_fd_sc_hd__or3_2 _23894_ (.A(_13411_),
    .B(_13693_),
    .C(_13695_),
    .X(_13696_));
 sky130_fd_sc_hd__o21ai_2 _23895_ (.A1(_13693_),
    .A2(_13695_),
    .B1(_13411_),
    .Y(_13697_));
 sky130_fd_sc_hd__inv_2 _23896_ (.A(_13456_),
    .Y(_13698_));
 sky130_fd_sc_hd__or2b_2 _23897_ (.A(_13425_),
    .B_N(_13424_),
    .X(_13699_));
 sky130_fd_sc_hd__and4_2 _23898_ (.A(iX[14]),
    .B(iX[15]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_13700_));
 sky130_fd_sc_hd__a22oi_2 _23899_ (.A1(iX[15]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[14]),
    .Y(_13701_));
 sky130_fd_sc_hd__nor2_2 _23900_ (.A(_13700_),
    .B(_13701_),
    .Y(_13702_));
 sky130_fd_sc_hd__nand2_2 _23901_ (.A(iX[13]),
    .B(iY[29]),
    .Y(_13703_));
 sky130_fd_sc_hd__xnor2_2 _23902_ (.A(_13702_),
    .B(_13703_),
    .Y(_13704_));
 sky130_fd_sc_hd__o21ba_2 _23903_ (.A1(_13421_),
    .A2(_13423_),
    .B1_N(_13419_),
    .X(_13706_));
 sky130_fd_sc_hd__xnor2_2 _23904_ (.A(_13704_),
    .B(_13706_),
    .Y(_13707_));
 sky130_fd_sc_hd__nand3_2 _23905_ (.A(iX[12]),
    .B(iY[30]),
    .C(_13707_),
    .Y(_13708_));
 sky130_fd_sc_hd__a21o_2 _23906_ (.A1(iX[12]),
    .A2(iY[30]),
    .B1(_13707_),
    .X(_13709_));
 sky130_fd_sc_hd__nand2_2 _23907_ (.A(_13708_),
    .B(_13709_),
    .Y(_13710_));
 sky130_fd_sc_hd__a21o_2 _23908_ (.A1(_13699_),
    .A2(_13427_),
    .B1(_13710_),
    .X(_13711_));
 sky130_fd_sc_hd__nand3_2 _23909_ (.A(_13699_),
    .B(_13427_),
    .C(_13710_),
    .Y(_13712_));
 sky130_fd_sc_hd__nand2_2 _23910_ (.A(_13711_),
    .B(_13712_),
    .Y(_13713_));
 sky130_fd_sc_hd__nand2_2 _23911_ (.A(iX[11]),
    .B(iY[31]),
    .Y(_13714_));
 sky130_fd_sc_hd__nand2_2 _23912_ (.A(_13713_),
    .B(_13714_),
    .Y(_13715_));
 sky130_fd_sc_hd__or2_2 _23913_ (.A(_13713_),
    .B(_13714_),
    .X(_13717_));
 sky130_fd_sc_hd__and2_2 _23914_ (.A(_13715_),
    .B(_13717_),
    .X(_13718_));
 sky130_fd_sc_hd__or2b_2 _23915_ (.A(_13441_),
    .B_N(_13447_),
    .X(_13719_));
 sky130_fd_sc_hd__or2b_2 _23916_ (.A(_13440_),
    .B_N(_13448_),
    .X(_13720_));
 sky130_fd_sc_hd__and2b_2 _23917_ (.A_N(_13384_),
    .B(_13383_),
    .X(_13721_));
 sky130_fd_sc_hd__o21ba_2 _23918_ (.A1(_13444_),
    .A2(_13446_),
    .B1_N(_13443_),
    .X(_13722_));
 sky130_fd_sc_hd__o21ba_2 _23919_ (.A1(_13374_),
    .A2(_13377_),
    .B1_N(_13373_),
    .X(_13723_));
 sky130_fd_sc_hd__and4_2 _23920_ (.A(iX[17]),
    .B(iX[18]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_13724_));
 sky130_fd_sc_hd__a22oi_2 _23921_ (.A1(iX[18]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[17]),
    .Y(_13725_));
 sky130_fd_sc_hd__nor2_2 _23922_ (.A(_13724_),
    .B(_13725_),
    .Y(_13726_));
 sky130_fd_sc_hd__nand2_2 _23923_ (.A(iX[16]),
    .B(iY[26]),
    .Y(_13728_));
 sky130_fd_sc_hd__xnor2_2 _23924_ (.A(_13726_),
    .B(_13728_),
    .Y(_13729_));
 sky130_fd_sc_hd__xnor2_2 _23925_ (.A(_13723_),
    .B(_13729_),
    .Y(_13730_));
 sky130_fd_sc_hd__xnor2_2 _23926_ (.A(_13722_),
    .B(_13730_),
    .Y(_13731_));
 sky130_fd_sc_hd__o21a_2 _23927_ (.A1(_13721_),
    .A2(_13386_),
    .B1(_13731_),
    .X(_13732_));
 sky130_fd_sc_hd__nor3_2 _23928_ (.A(_13721_),
    .B(_13386_),
    .C(_13731_),
    .Y(_13733_));
 sky130_fd_sc_hd__a211oi_2 _23929_ (.A1(_13719_),
    .A2(_13720_),
    .B1(_13732_),
    .C1(_13733_),
    .Y(_13734_));
 sky130_fd_sc_hd__o211a_2 _23930_ (.A1(_13732_),
    .A2(_13733_),
    .B1(_13719_),
    .C1(_13720_),
    .X(_13735_));
 sky130_fd_sc_hd__nor2_2 _23931_ (.A(_13450_),
    .B(_13452_),
    .Y(_13736_));
 sky130_fd_sc_hd__or3_2 _23932_ (.A(_13734_),
    .B(_13735_),
    .C(_13736_),
    .X(_13737_));
 sky130_fd_sc_hd__o21ai_2 _23933_ (.A1(_13734_),
    .A2(_13735_),
    .B1(_13736_),
    .Y(_13739_));
 sky130_fd_sc_hd__and3_2 _23934_ (.A(_13718_),
    .B(_13737_),
    .C(_13739_),
    .X(_13740_));
 sky130_fd_sc_hd__a21oi_2 _23935_ (.A1(_13737_),
    .A2(_13739_),
    .B1(_13718_),
    .Y(_13741_));
 sky130_fd_sc_hd__nor2_2 _23936_ (.A(_13740_),
    .B(_13741_),
    .Y(_13742_));
 sky130_fd_sc_hd__o21ai_2 _23937_ (.A1(_13406_),
    .A2(_13408_),
    .B1(_13742_),
    .Y(_13743_));
 sky130_fd_sc_hd__or3_2 _23938_ (.A(_13406_),
    .B(_13408_),
    .C(_13742_),
    .X(_13744_));
 sky130_fd_sc_hd__o211ai_2 _23939_ (.A1(_13698_),
    .A2(_13458_),
    .B1(_13743_),
    .C1(_13744_),
    .Y(_13745_));
 sky130_fd_sc_hd__a211o_2 _23940_ (.A1(_13743_),
    .A2(_13744_),
    .B1(_13698_),
    .C1(_13458_),
    .X(_13746_));
 sky130_fd_sc_hd__nand4_2 _23941_ (.A(_13696_),
    .B(_13697_),
    .C(_13745_),
    .D(_13746_),
    .Y(_13747_));
 sky130_fd_sc_hd__a22o_2 _23942_ (.A1(_13696_),
    .A2(_13697_),
    .B1(_13745_),
    .B2(_13746_),
    .X(_13748_));
 sky130_fd_sc_hd__nand2_2 _23943_ (.A(_13413_),
    .B(_13466_),
    .Y(_13750_));
 sky130_fd_sc_hd__and3_2 _23944_ (.A(_13747_),
    .B(_13748_),
    .C(_13750_),
    .X(_13751_));
 sky130_fd_sc_hd__a21oi_2 _23945_ (.A1(_13747_),
    .A2(_13748_),
    .B1(_13750_),
    .Y(_13752_));
 sky130_fd_sc_hd__a211oi_2 _23946_ (.A1(_13460_),
    .A2(_13463_),
    .B1(_13751_),
    .C1(_13752_),
    .Y(_13753_));
 sky130_fd_sc_hd__o211a_2 _23947_ (.A1(_13751_),
    .A2(_13752_),
    .B1(_13460_),
    .C1(_13463_),
    .X(_13754_));
 sky130_fd_sc_hd__nor2_2 _23948_ (.A(_13753_),
    .B(_13754_),
    .Y(_13755_));
 sky130_fd_sc_hd__o21ai_2 _23949_ (.A1(_13469_),
    .A2(_13471_),
    .B1(_13755_),
    .Y(_13756_));
 sky130_fd_sc_hd__or3_2 _23950_ (.A(_13469_),
    .B(_13471_),
    .C(_13755_),
    .X(_13757_));
 sky130_fd_sc_hd__and2_2 _23951_ (.A(_13756_),
    .B(_13757_),
    .X(_13758_));
 sky130_fd_sc_hd__o21ai_2 _23952_ (.A1(_13430_),
    .A2(_13435_),
    .B1(_13758_),
    .Y(_13759_));
 sky130_fd_sc_hd__or3_2 _23953_ (.A(_13430_),
    .B(_13435_),
    .C(_13758_),
    .X(_13761_));
 sky130_fd_sc_hd__nand2_2 _23954_ (.A(_13759_),
    .B(_13761_),
    .Y(_13762_));
 sky130_fd_sc_hd__o21bai_2 _23955_ (.A1(_13474_),
    .A2(_13479_),
    .B1_N(_13762_),
    .Y(_13763_));
 sky130_fd_sc_hd__or3b_2 _23956_ (.A(_13474_),
    .B(_13479_),
    .C_N(_13762_),
    .X(_13764_));
 sky130_fd_sc_hd__and2_2 _23957_ (.A(_13763_),
    .B(_13764_),
    .X(_13765_));
 sky130_fd_sc_hd__o21ba_2 _23958_ (.A1(_13481_),
    .A2(_13482_),
    .B1_N(_13484_),
    .X(_13766_));
 sky130_fd_sc_hd__o21ai_2 _23959_ (.A1(_13485_),
    .A2(_13483_),
    .B1(_13766_),
    .Y(_13767_));
 sky130_fd_sc_hd__xor2_2 _23960_ (.A(_13765_),
    .B(_13767_),
    .X(_13768_));
 sky130_fd_sc_hd__or2b_2 _23961_ (.A(_13613_),
    .B_N(_13612_),
    .X(_13769_));
 sky130_fd_sc_hd__nand2_2 _23962_ (.A(_13608_),
    .B(_13609_),
    .Y(_13770_));
 sky130_fd_sc_hd__nand2_2 _23963_ (.A(iY[33]),
    .B(iX[41]),
    .Y(_13772_));
 sky130_fd_sc_hd__a22o_2 _23964_ (.A1(iY[35]),
    .A2(iX[39]),
    .B1(iX[40]),
    .B2(iY[34]),
    .X(_13773_));
 sky130_fd_sc_hd__nand4_2 _23965_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[39]),
    .D(iX[40]),
    .Y(_13774_));
 sky130_fd_sc_hd__nand3b_2 _23966_ (.A_N(_13772_),
    .B(_13773_),
    .C(_13774_),
    .Y(_13775_));
 sky130_fd_sc_hd__a21bo_2 _23967_ (.A1(_13774_),
    .A2(_13773_),
    .B1_N(_13772_),
    .X(_13776_));
 sky130_fd_sc_hd__o21bai_2 _23968_ (.A1(_13568_),
    .A2(_13569_),
    .B1_N(_13567_),
    .Y(_13777_));
 sky130_fd_sc_hd__nand3_2 _23969_ (.A(_13775_),
    .B(_13776_),
    .C(_13777_),
    .Y(_13778_));
 sky130_fd_sc_hd__a21o_2 _23970_ (.A1(_13775_),
    .A2(_13776_),
    .B1(_13777_),
    .X(_13779_));
 sky130_fd_sc_hd__and4_2 _23971_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[38]),
    .D(iX[42]),
    .X(_13780_));
 sky130_fd_sc_hd__a22oi_2 _23972_ (.A1(iY[36]),
    .A2(iX[38]),
    .B1(iX[42]),
    .B2(iY[32]),
    .Y(_13781_));
 sky130_fd_sc_hd__or2_2 _23973_ (.A(_13780_),
    .B(_13781_),
    .X(_13783_));
 sky130_fd_sc_hd__nand2_2 _23974_ (.A(iX[37]),
    .B(iY[37]),
    .Y(_13784_));
 sky130_fd_sc_hd__xor2_2 _23975_ (.A(_13783_),
    .B(_13784_),
    .X(_13785_));
 sky130_fd_sc_hd__nand3_2 _23976_ (.A(_13778_),
    .B(_13779_),
    .C(_13785_),
    .Y(_13786_));
 sky130_fd_sc_hd__a21o_2 _23977_ (.A1(_13778_),
    .A2(_13779_),
    .B1(_13785_),
    .X(_13787_));
 sky130_fd_sc_hd__a21bo_2 _23978_ (.A1(_13575_),
    .A2(_13580_),
    .B1_N(_13573_),
    .X(_13788_));
 sky130_fd_sc_hd__nand3_2 _23979_ (.A(_13786_),
    .B(_13787_),
    .C(_13788_),
    .Y(_13789_));
 sky130_fd_sc_hd__a21o_2 _23980_ (.A1(_13786_),
    .A2(_13787_),
    .B1(_13788_),
    .X(_13790_));
 sky130_fd_sc_hd__o21ba_2 _23981_ (.A1(_13590_),
    .A2(_13592_),
    .B1_N(_13589_),
    .X(_13791_));
 sky130_fd_sc_hd__o21ba_2 _23982_ (.A1(_13577_),
    .A2(_13579_),
    .B1_N(_13576_),
    .X(_13792_));
 sky130_fd_sc_hd__and4_2 _23983_ (.A(iX[35]),
    .B(iX[36]),
    .C(iY[38]),
    .D(iY[39]),
    .X(_13794_));
 sky130_fd_sc_hd__a22oi_2 _23984_ (.A1(iX[36]),
    .A2(iY[38]),
    .B1(iY[39]),
    .B2(iX[35]),
    .Y(_13795_));
 sky130_fd_sc_hd__nor2_2 _23985_ (.A(_13794_),
    .B(_13795_),
    .Y(_13796_));
 sky130_fd_sc_hd__nand2_2 _23986_ (.A(iX[34]),
    .B(iY[40]),
    .Y(_13797_));
 sky130_fd_sc_hd__xnor2_2 _23987_ (.A(_13796_),
    .B(_13797_),
    .Y(_13798_));
 sky130_fd_sc_hd__xnor2_2 _23988_ (.A(_13792_),
    .B(_13798_),
    .Y(_13799_));
 sky130_fd_sc_hd__xnor2_2 _23989_ (.A(_13791_),
    .B(_13799_),
    .Y(_13800_));
 sky130_fd_sc_hd__and3_2 _23990_ (.A(_13789_),
    .B(_13790_),
    .C(_13800_),
    .X(_13801_));
 sky130_fd_sc_hd__a21oi_2 _23991_ (.A1(_13789_),
    .A2(_13790_),
    .B1(_13800_),
    .Y(_13802_));
 sky130_fd_sc_hd__a211o_2 _23992_ (.A1(_13584_),
    .A2(_13597_),
    .B1(_13801_),
    .C1(_13802_),
    .X(_13803_));
 sky130_fd_sc_hd__o211ai_2 _23993_ (.A1(_13801_),
    .A2(_13802_),
    .B1(_13584_),
    .C1(_13597_),
    .Y(_13805_));
 sky130_fd_sc_hd__or2b_2 _23994_ (.A(_13588_),
    .B_N(_13593_),
    .X(_13806_));
 sky130_fd_sc_hd__or2b_2 _23995_ (.A(_13587_),
    .B_N(_13594_),
    .X(_13807_));
 sky130_fd_sc_hd__a22oi_2 _23996_ (.A1(iX[33]),
    .A2(iY[41]),
    .B1(iY[42]),
    .B2(iX[32]),
    .Y(_13808_));
 sky130_fd_sc_hd__and4_2 _23997_ (.A(iX[33]),
    .B(iX[32]),
    .C(iY[41]),
    .D(iY[42]),
    .X(_13809_));
 sky130_fd_sc_hd__or2_2 _23998_ (.A(_13808_),
    .B(_13809_),
    .X(_13810_));
 sky130_fd_sc_hd__a21oi_2 _23999_ (.A1(_13806_),
    .A2(_13807_),
    .B1(_13810_),
    .Y(_13811_));
 sky130_fd_sc_hd__and3_2 _24000_ (.A(_13806_),
    .B(_13807_),
    .C(_13810_),
    .X(_13812_));
 sky130_fd_sc_hd__nor2_2 _24001_ (.A(_13811_),
    .B(_13812_),
    .Y(_13813_));
 sky130_fd_sc_hd__nand3_2 _24002_ (.A(_13803_),
    .B(_13805_),
    .C(_13813_),
    .Y(_13814_));
 sky130_fd_sc_hd__a21o_2 _24003_ (.A1(_13803_),
    .A2(_13805_),
    .B1(_13813_),
    .X(_13816_));
 sky130_fd_sc_hd__and2_2 _24004_ (.A(_13814_),
    .B(_13816_),
    .X(_13817_));
 sky130_fd_sc_hd__a21o_2 _24005_ (.A1(_13600_),
    .A2(_13606_),
    .B1(_13599_),
    .X(_13818_));
 sky130_fd_sc_hd__xnor2_2 _24006_ (.A(_13817_),
    .B(_13818_),
    .Y(_13819_));
 sky130_fd_sc_hd__xnor2_2 _24007_ (.A(_13604_),
    .B(_13819_),
    .Y(_13820_));
 sky130_fd_sc_hd__xor2_2 _24008_ (.A(_13770_),
    .B(_13820_),
    .X(_13821_));
 sky130_fd_sc_hd__or2_2 _24009_ (.A(_13566_),
    .B(_13610_),
    .X(_13822_));
 sky130_fd_sc_hd__nor2_2 _24010_ (.A(_13333_),
    .B(_13334_),
    .Y(_13823_));
 sky130_fd_sc_hd__or4b_2 _24011_ (.A(_12902_),
    .B(_13610_),
    .C(_13823_),
    .D_N(_13566_),
    .X(_13824_));
 sky130_fd_sc_hd__nand2_2 _24012_ (.A(_13822_),
    .B(_13824_),
    .Y(_13825_));
 sky130_fd_sc_hd__xor2_2 _24013_ (.A(_13821_),
    .B(_13825_),
    .X(_13827_));
 sky130_fd_sc_hd__xnor2_2 _24014_ (.A(_13769_),
    .B(_13827_),
    .Y(_13828_));
 sky130_fd_sc_hd__and2b_2 _24015_ (.A_N(_13337_),
    .B(_13297_),
    .X(_13829_));
 sky130_fd_sc_hd__a22oi_2 _24016_ (.A1(_13829_),
    .A2(_13612_),
    .B1(_13615_),
    .B2(_13339_),
    .Y(_13830_));
 sky130_fd_sc_hd__xnor2_2 _24017_ (.A(_13828_),
    .B(_13830_),
    .Y(_13831_));
 sky130_fd_sc_hd__nor3_2 _24018_ (.A(_13534_),
    .B(_13535_),
    .C(_13548_),
    .Y(_13832_));
 sky130_fd_sc_hd__nand3_2 _24019_ (.A(_13514_),
    .B(_13515_),
    .C(_13516_),
    .Y(_13833_));
 sky130_fd_sc_hd__or4_4 _24020_ (.A(_13517_),
    .B(_13518_),
    .C(_13529_),
    .D(_13531_),
    .X(_13834_));
 sky130_fd_sc_hd__and2_2 _24021_ (.A(iX[10]),
    .B(iX[42]),
    .X(_13835_));
 sky130_fd_sc_hd__nor2_2 _24022_ (.A(iX[10]),
    .B(iX[42]),
    .Y(_13836_));
 sky130_fd_sc_hd__nor2_2 _24023_ (.A(_13835_),
    .B(_13836_),
    .Y(_13838_));
 sky130_fd_sc_hd__nor3_2 _24024_ (.A(_13238_),
    .B(_13239_),
    .C(_13494_),
    .Y(_13839_));
 sky130_fd_sc_hd__o21ba_2 _24025_ (.A1(_13238_),
    .A2(_13491_),
    .B1_N(_13492_),
    .X(_13840_));
 sky130_fd_sc_hd__a21o_2 _24026_ (.A1(_13237_),
    .A2(_13839_),
    .B1(_13840_),
    .X(_13841_));
 sky130_fd_sc_hd__xnor2_2 _24027_ (.A(_13838_),
    .B(_13841_),
    .Y(_13842_));
 sky130_fd_sc_hd__or4_4 _24028_ (.A(_11565_),
    .B(_11574_),
    .C(_13502_),
    .D(_13842_),
    .X(_13843_));
 sky130_fd_sc_hd__xnor2_2 _24029_ (.A(iX[10]),
    .B(iX[42]),
    .Y(_13844_));
 sky130_fd_sc_hd__xnor2_2 _24030_ (.A(_13844_),
    .B(_13841_),
    .Y(_13845_));
 sky130_fd_sc_hd__a22o_2 _24031_ (.A1(_11582_),
    .A2(_13496_),
    .B1(_13845_),
    .B2(_11379_),
    .X(_13846_));
 sky130_fd_sc_hd__nand4_2 _24032_ (.A(_12451_),
    .B(_13244_),
    .C(_13843_),
    .D(_13846_),
    .Y(_13847_));
 sky130_fd_sc_hd__a22o_2 _24033_ (.A1(_12451_),
    .A2(_13244_),
    .B1(_13843_),
    .B2(_13846_),
    .X(_13849_));
 sky130_fd_sc_hd__a31o_2 _24034_ (.A1(_12451_),
    .A2(_13501_),
    .A3(_13499_),
    .B1(_13498_),
    .X(_13850_));
 sky130_fd_sc_hd__nand3_2 _24035_ (.A(_13847_),
    .B(_13849_),
    .C(_13850_),
    .Y(_13851_));
 sky130_fd_sc_hd__a21o_2 _24036_ (.A1(_13847_),
    .A2(_13849_),
    .B1(_13850_),
    .X(_13852_));
 sky130_fd_sc_hd__or4_2 _24037_ (.A(_12244_),
    .B(_12247_),
    .C(_13231_),
    .D(_12808_),
    .X(_13853_));
 sky130_fd_sc_hd__a22o_2 _24038_ (.A1(_12241_),
    .A2(_12810_),
    .B1(_13501_),
    .B2(_11842_),
    .X(_13854_));
 sky130_fd_sc_hd__nand2_2 _24039_ (.A(_13853_),
    .B(_13854_),
    .Y(_13855_));
 sky130_fd_sc_hd__nand2_2 _24040_ (.A(_12460_),
    .B(_12477_),
    .Y(_13856_));
 sky130_fd_sc_hd__xor2_2 _24041_ (.A(_13855_),
    .B(_13856_),
    .X(_13857_));
 sky130_fd_sc_hd__nand3_2 _24042_ (.A(_13851_),
    .B(_13852_),
    .C(_13857_),
    .Y(_13858_));
 sky130_fd_sc_hd__a21o_2 _24043_ (.A1(_13851_),
    .A2(_13852_),
    .B1(_13857_),
    .X(_13860_));
 sky130_fd_sc_hd__a21bo_2 _24044_ (.A1(_13507_),
    .A2(_13513_),
    .B1_N(_13506_),
    .X(_13861_));
 sky130_fd_sc_hd__and3_2 _24045_ (.A(_13858_),
    .B(_13860_),
    .C(_13861_),
    .X(_13862_));
 sky130_fd_sc_hd__a21oi_2 _24046_ (.A1(_13858_),
    .A2(_13860_),
    .B1(_13861_),
    .Y(_13863_));
 sky130_fd_sc_hd__or2b_2 _24047_ (.A(_13523_),
    .B_N(_13525_),
    .X(_13864_));
 sky130_fd_sc_hd__a31o_2 _24048_ (.A1(_12225_),
    .A2(_12759_),
    .A3(_13511_),
    .B1(_13509_),
    .X(_13865_));
 sky130_fd_sc_hd__nor2_2 _24049_ (.A(_12223_),
    .B(_12772_),
    .Y(_13866_));
 sky130_fd_sc_hd__or3b_2 _24050_ (.A(_11827_),
    .B(_12849_),
    .C_N(_13866_),
    .X(_13867_));
 sky130_fd_sc_hd__a21o_2 _24051_ (.A1(_11829_),
    .A2(_12845_),
    .B1(_13866_),
    .X(_13868_));
 sky130_fd_sc_hd__nand4_2 _24052_ (.A(_12827_),
    .B(_13274_),
    .C(_13867_),
    .D(_13868_),
    .Y(_13869_));
 sky130_fd_sc_hd__a22o_2 _24053_ (.A1(_11783_),
    .A2(_13274_),
    .B1(_13867_),
    .B2(_13868_),
    .X(_13871_));
 sky130_fd_sc_hd__nand3_2 _24054_ (.A(_13865_),
    .B(_13869_),
    .C(_13871_),
    .Y(_13872_));
 sky130_fd_sc_hd__a21o_2 _24055_ (.A1(_13869_),
    .A2(_13871_),
    .B1(_13865_),
    .X(_13873_));
 sky130_fd_sc_hd__and3_2 _24056_ (.A(_13864_),
    .B(_13872_),
    .C(_13873_),
    .X(_13874_));
 sky130_fd_sc_hd__a21oi_2 _24057_ (.A1(_13872_),
    .A2(_13873_),
    .B1(_13864_),
    .Y(_13875_));
 sky130_fd_sc_hd__nor4_2 _24058_ (.A(_13862_),
    .B(_13863_),
    .C(_13874_),
    .D(_13875_),
    .Y(_13876_));
 sky130_fd_sc_hd__o22a_2 _24059_ (.A1(_13862_),
    .A2(_13863_),
    .B1(_13874_),
    .B2(_13875_),
    .X(_13877_));
 sky130_fd_sc_hd__a211oi_2 _24060_ (.A1(_13833_),
    .A2(_13834_),
    .B1(_13876_),
    .C1(_13877_),
    .Y(_13878_));
 sky130_fd_sc_hd__o211a_2 _24061_ (.A1(_13876_),
    .A2(_13877_),
    .B1(_13833_),
    .C1(_13834_),
    .X(_13879_));
 sky130_fd_sc_hd__a21boi_2 _24062_ (.A1(_13520_),
    .A2(_13528_),
    .B1_N(_13527_),
    .Y(_13880_));
 sky130_fd_sc_hd__nand2_2 _24063_ (.A(iY[10]),
    .B(iY[42]),
    .Y(_13882_));
 sky130_fd_sc_hd__or2_2 _24064_ (.A(iY[10]),
    .B(iY[42]),
    .X(_13883_));
 sky130_fd_sc_hd__nand2_4 _24065_ (.A(_13882_),
    .B(_13883_),
    .Y(_13884_));
 sky130_fd_sc_hd__a22o_2 _24066_ (.A1(iY[8]),
    .A2(iY[40]),
    .B1(iY[41]),
    .B2(iY[9]),
    .X(_13885_));
 sky130_fd_sc_hd__o21a_2 _24067_ (.A1(_13539_),
    .A2(_13885_),
    .B1(_13536_),
    .X(_13886_));
 sky130_fd_sc_hd__xnor2_2 _24068_ (.A(_13884_),
    .B(_13886_),
    .Y(_13887_));
 sky130_fd_sc_hd__buf_1 _24069_ (.A(_13887_),
    .X(_13888_));
 sky130_fd_sc_hd__buf_1 _24070_ (.A(_13888_),
    .X(_13889_));
 sky130_fd_sc_hd__a22o_2 _24071_ (.A1(_12838_),
    .A2(_13544_),
    .B1(_13889_),
    .B2(_11374_),
    .X(_13890_));
 sky130_fd_sc_hd__xor2_2 _24072_ (.A(_13884_),
    .B(_13886_),
    .X(_13891_));
 sky130_fd_sc_hd__buf_1 _24073_ (.A(_13891_),
    .X(_13893_));
 sky130_fd_sc_hd__or3_2 _24074_ (.A(_11570_),
    .B(_13545_),
    .C(_13893_),
    .X(_13894_));
 sky130_fd_sc_hd__nand2_2 _24075_ (.A(_13890_),
    .B(_13894_),
    .Y(_13895_));
 sky130_fd_sc_hd__xnor2_2 _24076_ (.A(_13880_),
    .B(_13895_),
    .Y(_13896_));
 sky130_fd_sc_hd__or3_4 _24077_ (.A(_13878_),
    .B(_13879_),
    .C(_13896_),
    .X(_13897_));
 sky130_fd_sc_hd__o21ai_2 _24078_ (.A1(_13878_),
    .A2(_13879_),
    .B1(_13896_),
    .Y(_13898_));
 sky130_fd_sc_hd__o211ai_2 _24079_ (.A1(_13534_),
    .A2(_13832_),
    .B1(_13897_),
    .C1(_13898_),
    .Y(_13899_));
 sky130_fd_sc_hd__a211o_2 _24080_ (.A1(_13897_),
    .A2(_13898_),
    .B1(_13534_),
    .C1(_13832_),
    .X(_13900_));
 sky130_fd_sc_hd__nand3_2 _24081_ (.A(_13546_),
    .B(_13899_),
    .C(_13900_),
    .Y(_13901_));
 sky130_fd_sc_hd__a21o_2 _24082_ (.A1(_13899_),
    .A2(_13900_),
    .B1(_13546_),
    .X(_13902_));
 sky130_fd_sc_hd__and3_2 _24083_ (.A(_13551_),
    .B(_13901_),
    .C(_13902_),
    .X(_13904_));
 sky130_fd_sc_hd__a21o_2 _24084_ (.A1(_13901_),
    .A2(_13902_),
    .B1(_13551_),
    .X(_13905_));
 sky130_fd_sc_hd__nor2b_2 _24085_ (.A(_13904_),
    .B_N(_13905_),
    .Y(_13906_));
 sky130_fd_sc_hd__or2_2 _24086_ (.A(_13554_),
    .B(_13556_),
    .X(_13907_));
 sky130_fd_sc_hd__xnor2_2 _24087_ (.A(_13906_),
    .B(_13907_),
    .Y(_13908_));
 sky130_fd_sc_hd__a21boi_2 _24088_ (.A1(_13561_),
    .A2(_13560_),
    .B1_N(_13559_),
    .Y(_13909_));
 sky130_fd_sc_hd__and2_2 _24089_ (.A(_13908_),
    .B(_13909_),
    .X(_13910_));
 sky130_fd_sc_hd__nor2_2 _24090_ (.A(_13908_),
    .B(_13909_),
    .Y(_13911_));
 sky130_fd_sc_hd__nor2_2 _24091_ (.A(_13910_),
    .B(_13911_),
    .Y(_13912_));
 sky130_fd_sc_hd__xnor2_2 _24092_ (.A(_13831_),
    .B(_13912_),
    .Y(_13913_));
 sky130_fd_sc_hd__xor2_2 _24093_ (.A(oO[10]),
    .B(_13913_),
    .X(_13915_));
 sky130_fd_sc_hd__and2b_2 _24094_ (.A_N(_13617_),
    .B(_13620_),
    .X(_13916_));
 sky130_fd_sc_hd__xnor2_2 _24095_ (.A(_13915_),
    .B(_13916_),
    .Y(_13917_));
 sky130_fd_sc_hd__o21bai_2 _24096_ (.A1(_13625_),
    .A2(_13628_),
    .B1_N(_13624_),
    .Y(_13918_));
 sky130_fd_sc_hd__xor2_2 _24097_ (.A(_13917_),
    .B(_13918_),
    .X(_13919_));
 sky130_fd_sc_hd__nor2_2 _24098_ (.A(_13768_),
    .B(_13919_),
    .Y(_13920_));
 sky130_fd_sc_hd__and2_2 _24099_ (.A(_13768_),
    .B(_13919_),
    .X(_13921_));
 sky130_fd_sc_hd__nor2_2 _24100_ (.A(_13920_),
    .B(_13921_),
    .Y(_13922_));
 sky130_fd_sc_hd__xor2_2 _24101_ (.A(_13640_),
    .B(_13922_),
    .X(oO[42]));
 sky130_fd_sc_hd__nor2_2 _24102_ (.A(_13880_),
    .B(_13895_),
    .Y(_13923_));
 sky130_fd_sc_hd__a211o_2 _24103_ (.A1(_13833_),
    .A2(_13834_),
    .B1(_13876_),
    .C1(_13877_),
    .X(_13925_));
 sky130_fd_sc_hd__buf_1 _24104_ (.A(_12244_),
    .X(_13926_));
 sky130_fd_sc_hd__or4_2 _24105_ (.A(_13926_),
    .B(_12248_),
    .C(_12808_),
    .D(_13241_),
    .X(_13927_));
 sky130_fd_sc_hd__a22o_2 _24106_ (.A1(_12242_),
    .A2(_13501_),
    .B1(_13244_),
    .B2(_11842_),
    .X(_13928_));
 sky130_fd_sc_hd__nand2_2 _24107_ (.A(_13927_),
    .B(_13928_),
    .Y(_13929_));
 sky130_fd_sc_hd__nand2_2 _24108_ (.A(_12759_),
    .B(_12816_),
    .Y(_13930_));
 sky130_fd_sc_hd__xor2_2 _24109_ (.A(_13929_),
    .B(_13930_),
    .X(_13931_));
 sky130_fd_sc_hd__xnor2_2 _24110_ (.A(iX[11]),
    .B(iX[43]),
    .Y(_13932_));
 sky130_fd_sc_hd__a21oi_2 _24111_ (.A1(_13838_),
    .A2(_13841_),
    .B1(_13835_),
    .Y(_13933_));
 sky130_fd_sc_hd__xnor2_2 _24112_ (.A(_13932_),
    .B(_13933_),
    .Y(_13934_));
 sky130_fd_sc_hd__or4_2 _24113_ (.A(_11565_),
    .B(_11575_),
    .C(_13842_),
    .D(_13934_),
    .X(_13936_));
 sky130_fd_sc_hd__xor2_2 _24114_ (.A(_13932_),
    .B(_13933_),
    .X(_13937_));
 sky130_fd_sc_hd__buf_1 _24115_ (.A(_13937_),
    .X(_13938_));
 sky130_fd_sc_hd__a22o_2 _24116_ (.A1(_11583_),
    .A2(_13845_),
    .B1(_13938_),
    .B2(_11380_),
    .X(_13939_));
 sky130_fd_sc_hd__nand4_2 _24117_ (.A(_12451_),
    .B(_13496_),
    .C(_13936_),
    .D(_13939_),
    .Y(_13940_));
 sky130_fd_sc_hd__a22o_2 _24118_ (.A1(_12451_),
    .A2(_13496_),
    .B1(_13936_),
    .B2(_13939_),
    .X(_13941_));
 sky130_fd_sc_hd__nand2_2 _24119_ (.A(_13843_),
    .B(_13847_),
    .Y(_13942_));
 sky130_fd_sc_hd__nand3_2 _24120_ (.A(_13940_),
    .B(_13941_),
    .C(_13942_),
    .Y(_13943_));
 sky130_fd_sc_hd__a21o_2 _24121_ (.A1(_13940_),
    .A2(_13941_),
    .B1(_13942_),
    .X(_13944_));
 sky130_fd_sc_hd__nand3_2 _24122_ (.A(_13931_),
    .B(_13943_),
    .C(_13944_),
    .Y(_13945_));
 sky130_fd_sc_hd__a21o_2 _24123_ (.A1(_13943_),
    .A2(_13944_),
    .B1(_13931_),
    .X(_13947_));
 sky130_fd_sc_hd__nand2_2 _24124_ (.A(_13851_),
    .B(_13858_),
    .Y(_13948_));
 sky130_fd_sc_hd__nand3_2 _24125_ (.A(_13945_),
    .B(_13947_),
    .C(_13948_),
    .Y(_13949_));
 sky130_fd_sc_hd__a21o_2 _24126_ (.A1(_13945_),
    .A2(_13947_),
    .B1(_13948_),
    .X(_13950_));
 sky130_fd_sc_hd__nand2_2 _24127_ (.A(_13867_),
    .B(_13869_),
    .Y(_13951_));
 sky130_fd_sc_hd__o21ai_2 _24128_ (.A1(_13855_),
    .A2(_13856_),
    .B1(_13853_),
    .Y(_13952_));
 sky130_fd_sc_hd__nor2_2 _24129_ (.A(_12457_),
    .B(_12849_),
    .Y(_13953_));
 sky130_fd_sc_hd__o22a_2 _24130_ (.A1(_12457_),
    .A2(_12773_),
    .B1(_12850_),
    .B2(_12223_),
    .X(_13954_));
 sky130_fd_sc_hd__a21oi_2 _24131_ (.A1(_13866_),
    .A2(_13953_),
    .B1(_13954_),
    .Y(_13955_));
 sky130_fd_sc_hd__or2_2 _24132_ (.A(_11827_),
    .B(_13273_),
    .X(_13956_));
 sky130_fd_sc_hd__xnor2_2 _24133_ (.A(_13955_),
    .B(_13956_),
    .Y(_13958_));
 sky130_fd_sc_hd__xnor2_2 _24134_ (.A(_13952_),
    .B(_13958_),
    .Y(_13959_));
 sky130_fd_sc_hd__xnor2_2 _24135_ (.A(_13951_),
    .B(_13959_),
    .Y(_13960_));
 sky130_fd_sc_hd__nand3_2 _24136_ (.A(_13949_),
    .B(_13950_),
    .C(_13960_),
    .Y(_13961_));
 sky130_fd_sc_hd__a21o_2 _24137_ (.A1(_13949_),
    .A2(_13950_),
    .B1(_13960_),
    .X(_13962_));
 sky130_fd_sc_hd__or2_2 _24138_ (.A(_13862_),
    .B(_13876_),
    .X(_13963_));
 sky130_fd_sc_hd__and3_2 _24139_ (.A(_13961_),
    .B(_13962_),
    .C(_13963_),
    .X(_13964_));
 sky130_fd_sc_hd__a21oi_2 _24140_ (.A1(_13961_),
    .A2(_13962_),
    .B1(_13963_),
    .Y(_13965_));
 sky130_fd_sc_hd__and3_2 _24141_ (.A(_13865_),
    .B(_13869_),
    .C(_13871_),
    .X(_13966_));
 sky130_fd_sc_hd__and4_2 _24142_ (.A(_11581_),
    .B(_12827_),
    .C(_13542_),
    .D(_13887_),
    .X(_13967_));
 sky130_fd_sc_hd__a22o_2 _24143_ (.A1(_12827_),
    .A2(_13542_),
    .B1(_13888_),
    .B2(_11581_),
    .X(_13968_));
 sky130_fd_sc_hd__and2b_2 _24144_ (.A_N(_13967_),
    .B(_13968_),
    .X(_13969_));
 sky130_fd_sc_hd__xnor2_2 _24145_ (.A(iY[11]),
    .B(iY[43]),
    .Y(_13970_));
 sky130_fd_sc_hd__a21bo_2 _24146_ (.A1(_13883_),
    .A2(_13886_),
    .B1_N(_13882_),
    .X(_13971_));
 sky130_fd_sc_hd__xor2_2 _24147_ (.A(_13970_),
    .B(_13971_),
    .X(_13972_));
 sky130_fd_sc_hd__nor2_2 _24148_ (.A(_11577_),
    .B(_13972_),
    .Y(_13973_));
 sky130_fd_sc_hd__xnor2_2 _24149_ (.A(_13969_),
    .B(_13973_),
    .Y(_13974_));
 sky130_fd_sc_hd__xor2_2 _24150_ (.A(_13894_),
    .B(_13974_),
    .X(_13975_));
 sky130_fd_sc_hd__o21a_2 _24151_ (.A1(_13966_),
    .A2(_13874_),
    .B1(_13975_),
    .X(_13976_));
 sky130_fd_sc_hd__nor3_2 _24152_ (.A(_13966_),
    .B(_13874_),
    .C(_13975_),
    .Y(_13977_));
 sky130_fd_sc_hd__or2_2 _24153_ (.A(_13976_),
    .B(_13977_),
    .X(_13979_));
 sky130_fd_sc_hd__nor3_2 _24154_ (.A(_13964_),
    .B(_13965_),
    .C(_13979_),
    .Y(_13980_));
 sky130_fd_sc_hd__o21a_2 _24155_ (.A1(_13964_),
    .A2(_13965_),
    .B1(_13979_),
    .X(_13981_));
 sky130_fd_sc_hd__a211o_2 _24156_ (.A1(_13925_),
    .A2(_13897_),
    .B1(_13980_),
    .C1(_13981_),
    .X(_13982_));
 sky130_fd_sc_hd__o211ai_2 _24157_ (.A1(_13980_),
    .A2(_13981_),
    .B1(_13925_),
    .C1(_13897_),
    .Y(_13983_));
 sky130_fd_sc_hd__and3_2 _24158_ (.A(_13923_),
    .B(_13982_),
    .C(_13983_),
    .X(_13984_));
 sky130_fd_sc_hd__a21oi_2 _24159_ (.A1(_13982_),
    .A2(_13983_),
    .B1(_13923_),
    .Y(_13985_));
 sky130_fd_sc_hd__nand2_2 _24160_ (.A(_13899_),
    .B(_13901_),
    .Y(_13986_));
 sky130_fd_sc_hd__nor3b_2 _24161_ (.A(_13984_),
    .B(_13985_),
    .C_N(_13986_),
    .Y(_13987_));
 sky130_fd_sc_hd__o21ba_2 _24162_ (.A1(_13984_),
    .A2(_13985_),
    .B1_N(_13986_),
    .X(_13988_));
 sky130_fd_sc_hd__a21o_2 _24163_ (.A1(_13554_),
    .A2(_13905_),
    .B1(_13904_),
    .X(_13990_));
 sky130_fd_sc_hd__or3_2 _24164_ (.A(_13987_),
    .B(_13988_),
    .C(_13990_),
    .X(_13991_));
 sky130_fd_sc_hd__o21ai_2 _24165_ (.A1(_13987_),
    .A2(_13988_),
    .B1(_13990_),
    .Y(_13992_));
 sky130_fd_sc_hd__nand2_2 _24166_ (.A(_13556_),
    .B(_13906_),
    .Y(_13993_));
 sky130_fd_sc_hd__a21oi_2 _24167_ (.A1(_13991_),
    .A2(_13992_),
    .B1(_13993_),
    .Y(_13994_));
 sky130_fd_sc_hd__and3_2 _24168_ (.A(_13993_),
    .B(_13991_),
    .C(_13992_),
    .X(_13995_));
 sky130_fd_sc_hd__o21bai_2 _24169_ (.A1(_13994_),
    .A2(_13995_),
    .B1_N(_13911_),
    .Y(_13996_));
 sky130_fd_sc_hd__or3b_4 _24170_ (.A(_13994_),
    .B(_13995_),
    .C_N(_13911_),
    .X(_13997_));
 sky130_fd_sc_hd__or2_2 _24171_ (.A(_13824_),
    .B(_13821_),
    .X(_13998_));
 sky130_fd_sc_hd__and4_2 _24172_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[40]),
    .D(iX[41]),
    .X(_13999_));
 sky130_fd_sc_hd__a22oi_2 _24173_ (.A1(iY[35]),
    .A2(iX[40]),
    .B1(iX[41]),
    .B2(iY[34]),
    .Y(_14001_));
 sky130_fd_sc_hd__nor2_2 _24174_ (.A(_13999_),
    .B(_14001_),
    .Y(_14002_));
 sky130_fd_sc_hd__nand2_2 _24175_ (.A(iY[33]),
    .B(iX[42]),
    .Y(_14003_));
 sky130_fd_sc_hd__xnor2_2 _24176_ (.A(_14002_),
    .B(_14003_),
    .Y(_14004_));
 sky130_fd_sc_hd__nand2_2 _24177_ (.A(_13774_),
    .B(_13775_),
    .Y(_14005_));
 sky130_fd_sc_hd__xor2_2 _24178_ (.A(_14004_),
    .B(_14005_),
    .X(_14006_));
 sky130_fd_sc_hd__and4_2 _24179_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[39]),
    .D(iX[43]),
    .X(_14007_));
 sky130_fd_sc_hd__a22oi_2 _24180_ (.A1(iY[36]),
    .A2(iX[39]),
    .B1(iX[43]),
    .B2(iY[32]),
    .Y(_14008_));
 sky130_fd_sc_hd__nor2_2 _24181_ (.A(_14007_),
    .B(_14008_),
    .Y(_14009_));
 sky130_fd_sc_hd__nand2_2 _24182_ (.A(iY[37]),
    .B(iX[38]),
    .Y(_14010_));
 sky130_fd_sc_hd__xnor2_2 _24183_ (.A(_14009_),
    .B(_14010_),
    .Y(_14012_));
 sky130_fd_sc_hd__xnor2_2 _24184_ (.A(_14006_),
    .B(_14012_),
    .Y(_14013_));
 sky130_fd_sc_hd__a21o_2 _24185_ (.A1(_13778_),
    .A2(_13786_),
    .B1(_14013_),
    .X(_14014_));
 sky130_fd_sc_hd__nand3_2 _24186_ (.A(_13778_),
    .B(_13786_),
    .C(_14013_),
    .Y(_14015_));
 sky130_fd_sc_hd__o21ba_2 _24187_ (.A1(_13795_),
    .A2(_13797_),
    .B1_N(_13794_),
    .X(_14016_));
 sky130_fd_sc_hd__nor2_2 _24188_ (.A(_13783_),
    .B(_13784_),
    .Y(_14017_));
 sky130_fd_sc_hd__and4_2 _24189_ (.A(iX[36]),
    .B(iX[37]),
    .C(iY[38]),
    .D(iY[39]),
    .X(_14018_));
 sky130_fd_sc_hd__a22oi_2 _24190_ (.A1(iX[37]),
    .A2(iY[38]),
    .B1(iY[39]),
    .B2(iX[36]),
    .Y(_14019_));
 sky130_fd_sc_hd__nor2_2 _24191_ (.A(_14018_),
    .B(_14019_),
    .Y(_14020_));
 sky130_fd_sc_hd__nand2_2 _24192_ (.A(iX[35]),
    .B(iY[40]),
    .Y(_14021_));
 sky130_fd_sc_hd__xnor2_2 _24193_ (.A(_14020_),
    .B(_14021_),
    .Y(_14023_));
 sky130_fd_sc_hd__o21ai_2 _24194_ (.A1(_13780_),
    .A2(_14017_),
    .B1(_14023_),
    .Y(_14024_));
 sky130_fd_sc_hd__or3_2 _24195_ (.A(_13780_),
    .B(_14017_),
    .C(_14023_),
    .X(_14025_));
 sky130_fd_sc_hd__and2_2 _24196_ (.A(_14024_),
    .B(_14025_),
    .X(_14026_));
 sky130_fd_sc_hd__xnor2_2 _24197_ (.A(_14016_),
    .B(_14026_),
    .Y(_14027_));
 sky130_fd_sc_hd__nand3_2 _24198_ (.A(_14014_),
    .B(_14015_),
    .C(_14027_),
    .Y(_14028_));
 sky130_fd_sc_hd__a21o_2 _24199_ (.A1(_14014_),
    .A2(_14015_),
    .B1(_14027_),
    .X(_14029_));
 sky130_fd_sc_hd__a31o_2 _24200_ (.A1(_13786_),
    .A2(_13787_),
    .A3(_13788_),
    .B1(_13801_),
    .X(_14030_));
 sky130_fd_sc_hd__nand3_2 _24201_ (.A(_14028_),
    .B(_14029_),
    .C(_14030_),
    .Y(_14031_));
 sky130_fd_sc_hd__a21o_2 _24202_ (.A1(_14028_),
    .A2(_14029_),
    .B1(_14030_),
    .X(_14032_));
 sky130_fd_sc_hd__or2b_2 _24203_ (.A(_13792_),
    .B_N(_13798_),
    .X(_14034_));
 sky130_fd_sc_hd__or2b_2 _24204_ (.A(_13791_),
    .B_N(_13799_),
    .X(_14035_));
 sky130_fd_sc_hd__and4_2 _24205_ (.A(iX[33]),
    .B(iX[34]),
    .C(iY[41]),
    .D(iY[42]),
    .X(_14036_));
 sky130_fd_sc_hd__a22oi_2 _24206_ (.A1(iX[34]),
    .A2(iY[41]),
    .B1(iY[42]),
    .B2(iX[33]),
    .Y(_14037_));
 sky130_fd_sc_hd__nor2_2 _24207_ (.A(_14036_),
    .B(_14037_),
    .Y(_14038_));
 sky130_fd_sc_hd__nand2_2 _24208_ (.A(iX[32]),
    .B(iY[43]),
    .Y(_14039_));
 sky130_fd_sc_hd__xnor2_2 _24209_ (.A(_14038_),
    .B(_14039_),
    .Y(_14040_));
 sky130_fd_sc_hd__and2_2 _24210_ (.A(_13809_),
    .B(_14040_),
    .X(_14041_));
 sky130_fd_sc_hd__nor2_2 _24211_ (.A(_13809_),
    .B(_14040_),
    .Y(_14042_));
 sky130_fd_sc_hd__or2_2 _24212_ (.A(_14041_),
    .B(_14042_),
    .X(_14043_));
 sky130_fd_sc_hd__a21oi_2 _24213_ (.A1(_14034_),
    .A2(_14035_),
    .B1(_14043_),
    .Y(_14045_));
 sky130_fd_sc_hd__and3_2 _24214_ (.A(_14034_),
    .B(_14035_),
    .C(_14043_),
    .X(_14046_));
 sky130_fd_sc_hd__nor2_2 _24215_ (.A(_14045_),
    .B(_14046_),
    .Y(_14047_));
 sky130_fd_sc_hd__nand3_2 _24216_ (.A(_14031_),
    .B(_14032_),
    .C(_14047_),
    .Y(_14048_));
 sky130_fd_sc_hd__a21o_2 _24217_ (.A1(_14031_),
    .A2(_14032_),
    .B1(_14047_),
    .X(_14049_));
 sky130_fd_sc_hd__nand2_2 _24218_ (.A(_13803_),
    .B(_13814_),
    .Y(_14050_));
 sky130_fd_sc_hd__nand3_2 _24219_ (.A(_14048_),
    .B(_14049_),
    .C(_14050_),
    .Y(_14051_));
 sky130_fd_sc_hd__a21o_2 _24220_ (.A1(_14048_),
    .A2(_14049_),
    .B1(_14050_),
    .X(_14052_));
 sky130_fd_sc_hd__a21o_2 _24221_ (.A1(_14051_),
    .A2(_14052_),
    .B1(_13811_),
    .X(_14053_));
 sky130_fd_sc_hd__nand3_2 _24222_ (.A(_13811_),
    .B(_14051_),
    .C(_14052_),
    .Y(_14054_));
 sky130_fd_sc_hd__and2_2 _24223_ (.A(_14053_),
    .B(_14054_),
    .X(_14056_));
 sky130_fd_sc_hd__or2_2 _24224_ (.A(_13817_),
    .B(_13818_),
    .X(_14057_));
 sky130_fd_sc_hd__and3_2 _24225_ (.A(_13814_),
    .B(_13816_),
    .C(_13818_),
    .X(_14058_));
 sky130_fd_sc_hd__a21o_2 _24226_ (.A1(_13604_),
    .A2(_14057_),
    .B1(_14058_),
    .X(_14059_));
 sky130_fd_sc_hd__xnor2_2 _24227_ (.A(_14056_),
    .B(_14059_),
    .Y(_14060_));
 sky130_fd_sc_hd__or2b_2 _24228_ (.A(_13770_),
    .B_N(_13820_),
    .X(_14061_));
 sky130_fd_sc_hd__o21a_2 _24229_ (.A1(_13822_),
    .A2(_13821_),
    .B1(_14061_),
    .X(_14062_));
 sky130_fd_sc_hd__xnor2_2 _24230_ (.A(_14060_),
    .B(_14062_),
    .Y(_14063_));
 sky130_fd_sc_hd__or2_2 _24231_ (.A(_13998_),
    .B(_14063_),
    .X(_14064_));
 sky130_fd_sc_hd__nand2_2 _24232_ (.A(_13998_),
    .B(_14063_),
    .Y(_14065_));
 sky130_fd_sc_hd__nand2_2 _24233_ (.A(_14064_),
    .B(_14065_),
    .Y(_14067_));
 sky130_fd_sc_hd__or2_2 _24234_ (.A(_13769_),
    .B(_13827_),
    .X(_14068_));
 sky130_fd_sc_hd__o21ai_2 _24235_ (.A1(_13828_),
    .A2(_13830_),
    .B1(_14068_),
    .Y(_14069_));
 sky130_fd_sc_hd__xor2_2 _24236_ (.A(_14067_),
    .B(_14069_),
    .X(_14070_));
 sky130_fd_sc_hd__and3_2 _24237_ (.A(_13996_),
    .B(_13997_),
    .C(_14070_),
    .X(_14071_));
 sky130_fd_sc_hd__a21oi_2 _24238_ (.A1(_13996_),
    .A2(_13997_),
    .B1(_14070_),
    .Y(_14072_));
 sky130_fd_sc_hd__or2_2 _24239_ (.A(_14071_),
    .B(_14072_),
    .X(_14073_));
 sky130_fd_sc_hd__xnor2_2 _24240_ (.A(oO[11]),
    .B(_14073_),
    .Y(_14074_));
 sky130_fd_sc_hd__nand2_2 _24241_ (.A(_13831_),
    .B(_13912_),
    .Y(_14075_));
 sky130_fd_sc_hd__o21ai_2 _24242_ (.A1(oO[10]),
    .A2(_13913_),
    .B1(_14075_),
    .Y(_14076_));
 sky130_fd_sc_hd__xor2_2 _24243_ (.A(_14074_),
    .B(_14076_),
    .X(_14078_));
 sky130_fd_sc_hd__or2b_2 _24244_ (.A(_13916_),
    .B_N(_13915_),
    .X(_14079_));
 sky130_fd_sc_hd__a21boi_2 _24245_ (.A1(_13917_),
    .A2(_13918_),
    .B1_N(_14079_),
    .Y(_14080_));
 sky130_fd_sc_hd__nor2_2 _24246_ (.A(_14078_),
    .B(_14080_),
    .Y(_14081_));
 sky130_fd_sc_hd__and2_2 _24247_ (.A(_14078_),
    .B(_14080_),
    .X(_14082_));
 sky130_fd_sc_hd__a21oi_2 _24248_ (.A1(_13642_),
    .A2(_13648_),
    .B1(_13353_),
    .Y(_14083_));
 sky130_fd_sc_hd__and3_2 _24249_ (.A(iY[12]),
    .B(iX[31]),
    .C(_13643_),
    .X(_14084_));
 sky130_fd_sc_hd__a21oi_2 _24250_ (.A1(iY[12]),
    .A2(iX[31]),
    .B1(_13643_),
    .Y(_14085_));
 sky130_fd_sc_hd__and4bb_2 _24251_ (.A_N(_14084_),
    .B_N(_14085_),
    .C(iY[14]),
    .D(iX[29]),
    .X(_14086_));
 sky130_fd_sc_hd__o2bb2a_2 _24252_ (.A1_N(iY[14]),
    .A2_N(iX[29]),
    .B1(_14084_),
    .B2(_14085_),
    .X(_14087_));
 sky130_fd_sc_hd__nor2_2 _24253_ (.A(_14086_),
    .B(_14087_),
    .Y(_14089_));
 sky130_fd_sc_hd__and2b_2 _24254_ (.A_N(_14083_),
    .B(_14089_),
    .X(_14090_));
 sky130_fd_sc_hd__and2b_2 _24255_ (.A_N(_14089_),
    .B(_14083_),
    .X(_14091_));
 sky130_fd_sc_hd__nor2_2 _24256_ (.A(_14090_),
    .B(_14091_),
    .Y(_14092_));
 sky130_fd_sc_hd__a21o_2 _24257_ (.A1(_13397_),
    .A2(_13671_),
    .B1(_13682_),
    .X(_14093_));
 sky130_fd_sc_hd__and4_2 _24258_ (.A(iX[21]),
    .B(iY[21]),
    .C(iX[22]),
    .D(iY[22]),
    .X(_14094_));
 sky130_fd_sc_hd__a22oi_2 _24259_ (.A1(iY[21]),
    .A2(iX[22]),
    .B1(iY[22]),
    .B2(iX[21]),
    .Y(_14095_));
 sky130_fd_sc_hd__nor2_2 _24260_ (.A(_14094_),
    .B(_14095_),
    .Y(_14096_));
 sky130_fd_sc_hd__nand2_2 _24261_ (.A(iX[20]),
    .B(iY[23]),
    .Y(_14097_));
 sky130_fd_sc_hd__xnor2_2 _24262_ (.A(_14096_),
    .B(_14097_),
    .Y(_14098_));
 sky130_fd_sc_hd__and4_2 _24263_ (.A(iY[18]),
    .B(iY[19]),
    .C(iX[24]),
    .D(iX[25]),
    .X(_14100_));
 sky130_fd_sc_hd__a22oi_2 _24264_ (.A1(iY[19]),
    .A2(iX[24]),
    .B1(iX[25]),
    .B2(iY[18]),
    .Y(_14101_));
 sky130_fd_sc_hd__nor2_2 _24265_ (.A(_14100_),
    .B(_14101_),
    .Y(_14102_));
 sky130_fd_sc_hd__nand2_2 _24266_ (.A(iY[20]),
    .B(iX[23]),
    .Y(_14103_));
 sky130_fd_sc_hd__xnor2_2 _24267_ (.A(_14102_),
    .B(_14103_),
    .Y(_14104_));
 sky130_fd_sc_hd__o21ba_2 _24268_ (.A1(_13662_),
    .A2(_13664_),
    .B1_N(_13660_),
    .X(_14105_));
 sky130_fd_sc_hd__xnor2_2 _24269_ (.A(_14104_),
    .B(_14105_),
    .Y(_14106_));
 sky130_fd_sc_hd__and2_2 _24270_ (.A(_14098_),
    .B(_14106_),
    .X(_14107_));
 sky130_fd_sc_hd__nor2_2 _24271_ (.A(_14098_),
    .B(_14106_),
    .Y(_14108_));
 sky130_fd_sc_hd__or2_2 _24272_ (.A(_14107_),
    .B(_14108_),
    .X(_14109_));
 sky130_fd_sc_hd__or2b_2 _24273_ (.A(_13673_),
    .B_N(_13678_),
    .X(_14111_));
 sky130_fd_sc_hd__a31o_2 _24274_ (.A1(iY[17]),
    .A2(iX[25]),
    .A3(_13676_),
    .B1(_13674_),
    .X(_14112_));
 sky130_fd_sc_hd__and4_2 _24275_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[27]),
    .D(iX[28]),
    .X(_14113_));
 sky130_fd_sc_hd__a22oi_2 _24276_ (.A1(iY[16]),
    .A2(iX[27]),
    .B1(iX[28]),
    .B2(iY[15]),
    .Y(_14114_));
 sky130_fd_sc_hd__nor2_2 _24277_ (.A(_14113_),
    .B(_14114_),
    .Y(_14115_));
 sky130_fd_sc_hd__nand2_2 _24278_ (.A(iY[17]),
    .B(iX[26]),
    .Y(_14116_));
 sky130_fd_sc_hd__xnor2_2 _24279_ (.A(_14115_),
    .B(_14116_),
    .Y(_14117_));
 sky130_fd_sc_hd__o21ai_2 _24280_ (.A1(_13644_),
    .A2(_13646_),
    .B1(_14117_),
    .Y(_14118_));
 sky130_fd_sc_hd__or3_2 _24281_ (.A(_13644_),
    .B(_13646_),
    .C(_14117_),
    .X(_14119_));
 sky130_fd_sc_hd__and2_2 _24282_ (.A(_14118_),
    .B(_14119_),
    .X(_14120_));
 sky130_fd_sc_hd__xnor2_2 _24283_ (.A(_14112_),
    .B(_14120_),
    .Y(_14122_));
 sky130_fd_sc_hd__a21oi_2 _24284_ (.A1(_14111_),
    .A2(_13680_),
    .B1(_14122_),
    .Y(_14123_));
 sky130_fd_sc_hd__and3_2 _24285_ (.A(_14111_),
    .B(_13680_),
    .C(_14122_),
    .X(_14124_));
 sky130_fd_sc_hd__or3_2 _24286_ (.A(_14109_),
    .B(_14123_),
    .C(_14124_),
    .X(_14125_));
 sky130_fd_sc_hd__o21ai_2 _24287_ (.A1(_14123_),
    .A2(_14124_),
    .B1(_14109_),
    .Y(_14126_));
 sky130_fd_sc_hd__and3_2 _24288_ (.A(_13651_),
    .B(_14125_),
    .C(_14126_),
    .X(_14127_));
 sky130_fd_sc_hd__a21oi_2 _24289_ (.A1(_14125_),
    .A2(_14126_),
    .B1(_13651_),
    .Y(_14128_));
 sky130_fd_sc_hd__a211o_2 _24290_ (.A1(_14093_),
    .A2(_13686_),
    .B1(_14127_),
    .C1(_14128_),
    .X(_14129_));
 sky130_fd_sc_hd__o211ai_2 _24291_ (.A1(_14127_),
    .A2(_14128_),
    .B1(_14093_),
    .C1(_13686_),
    .Y(_14130_));
 sky130_fd_sc_hd__and3_2 _24292_ (.A(_14092_),
    .B(_14129_),
    .C(_14130_),
    .X(_14131_));
 sky130_fd_sc_hd__a21oi_2 _24293_ (.A1(_14129_),
    .A2(_14130_),
    .B1(_14092_),
    .Y(_14133_));
 sky130_fd_sc_hd__or3_2 _24294_ (.A(_13692_),
    .B(_14131_),
    .C(_14133_),
    .X(_14134_));
 sky130_fd_sc_hd__o21ai_2 _24295_ (.A1(_14131_),
    .A2(_14133_),
    .B1(_13692_),
    .Y(_14135_));
 sky130_fd_sc_hd__inv_2 _24296_ (.A(_13737_),
    .Y(_14136_));
 sky130_fd_sc_hd__or2b_2 _24297_ (.A(_13706_),
    .B_N(_13704_),
    .X(_14137_));
 sky130_fd_sc_hd__and4_2 _24298_ (.A(iX[15]),
    .B(iX[16]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_14138_));
 sky130_fd_sc_hd__a22oi_2 _24299_ (.A1(iX[16]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[15]),
    .Y(_14139_));
 sky130_fd_sc_hd__nor2_2 _24300_ (.A(_14138_),
    .B(_14139_),
    .Y(_14140_));
 sky130_fd_sc_hd__nand2_2 _24301_ (.A(iX[14]),
    .B(iY[29]),
    .Y(_14141_));
 sky130_fd_sc_hd__xnor2_2 _24302_ (.A(_14140_),
    .B(_14141_),
    .Y(_14142_));
 sky130_fd_sc_hd__o21ba_2 _24303_ (.A1(_13701_),
    .A2(_13703_),
    .B1_N(_13700_),
    .X(_14144_));
 sky130_fd_sc_hd__xnor2_2 _24304_ (.A(_14142_),
    .B(_14144_),
    .Y(_14145_));
 sky130_fd_sc_hd__nand3_2 _24305_ (.A(iX[13]),
    .B(iY[30]),
    .C(_14145_),
    .Y(_14146_));
 sky130_fd_sc_hd__a21o_2 _24306_ (.A1(iX[13]),
    .A2(iY[30]),
    .B1(_14145_),
    .X(_14147_));
 sky130_fd_sc_hd__nand2_2 _24307_ (.A(_14146_),
    .B(_14147_),
    .Y(_14148_));
 sky130_fd_sc_hd__a21oi_2 _24308_ (.A1(_14137_),
    .A2(_13708_),
    .B1(_14148_),
    .Y(_14149_));
 sky130_fd_sc_hd__and3_2 _24309_ (.A(_14137_),
    .B(_13708_),
    .C(_14148_),
    .X(_14150_));
 sky130_fd_sc_hd__nor2_2 _24310_ (.A(_14149_),
    .B(_14150_),
    .Y(_14151_));
 sky130_fd_sc_hd__a21oi_2 _24311_ (.A1(iX[12]),
    .A2(iY[31]),
    .B1(_14151_),
    .Y(_14152_));
 sky130_fd_sc_hd__and3_2 _24312_ (.A(iX[12]),
    .B(iY[31]),
    .C(_14151_),
    .X(_14153_));
 sky130_fd_sc_hd__nor2_2 _24313_ (.A(_14152_),
    .B(_14153_),
    .Y(_14155_));
 sky130_fd_sc_hd__or2b_2 _24314_ (.A(_13723_),
    .B_N(_13729_),
    .X(_14156_));
 sky130_fd_sc_hd__or2b_2 _24315_ (.A(_13722_),
    .B_N(_13730_),
    .X(_14157_));
 sky130_fd_sc_hd__and2b_2 _24316_ (.A_N(_13666_),
    .B(_13665_),
    .X(_14158_));
 sky130_fd_sc_hd__o21ba_2 _24317_ (.A1(_13725_),
    .A2(_13728_),
    .B1_N(_13724_),
    .X(_14159_));
 sky130_fd_sc_hd__o21ba_2 _24318_ (.A1(_13656_),
    .A2(_13658_),
    .B1_N(_13655_),
    .X(_14160_));
 sky130_fd_sc_hd__and4_2 _24319_ (.A(iX[18]),
    .B(iX[19]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_14161_));
 sky130_fd_sc_hd__a22oi_2 _24320_ (.A1(iX[19]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[18]),
    .Y(_14162_));
 sky130_fd_sc_hd__nor2_2 _24321_ (.A(_14161_),
    .B(_14162_),
    .Y(_14163_));
 sky130_fd_sc_hd__nand2_2 _24322_ (.A(iX[17]),
    .B(iY[26]),
    .Y(_14164_));
 sky130_fd_sc_hd__xnor2_2 _24323_ (.A(_14163_),
    .B(_14164_),
    .Y(_14166_));
 sky130_fd_sc_hd__xnor2_2 _24324_ (.A(_14160_),
    .B(_14166_),
    .Y(_14167_));
 sky130_fd_sc_hd__xnor2_2 _24325_ (.A(_14159_),
    .B(_14167_),
    .Y(_14168_));
 sky130_fd_sc_hd__o21a_2 _24326_ (.A1(_14158_),
    .A2(_13668_),
    .B1(_14168_),
    .X(_14169_));
 sky130_fd_sc_hd__nor3_2 _24327_ (.A(_14158_),
    .B(_13668_),
    .C(_14168_),
    .Y(_14170_));
 sky130_fd_sc_hd__a211oi_2 _24328_ (.A1(_14156_),
    .A2(_14157_),
    .B1(_14169_),
    .C1(_14170_),
    .Y(_14171_));
 sky130_fd_sc_hd__o211a_2 _24329_ (.A1(_14169_),
    .A2(_14170_),
    .B1(_14156_),
    .C1(_14157_),
    .X(_14172_));
 sky130_fd_sc_hd__nor2_2 _24330_ (.A(_13732_),
    .B(_13734_),
    .Y(_14173_));
 sky130_fd_sc_hd__or3_2 _24331_ (.A(_14171_),
    .B(_14172_),
    .C(_14173_),
    .X(_14174_));
 sky130_fd_sc_hd__o21ai_2 _24332_ (.A1(_14171_),
    .A2(_14172_),
    .B1(_14173_),
    .Y(_14175_));
 sky130_fd_sc_hd__and3_2 _24333_ (.A(_14155_),
    .B(_14174_),
    .C(_14175_),
    .X(_14177_));
 sky130_fd_sc_hd__a21oi_2 _24334_ (.A1(_14174_),
    .A2(_14175_),
    .B1(_14155_),
    .Y(_14178_));
 sky130_fd_sc_hd__nor2_2 _24335_ (.A(_14177_),
    .B(_14178_),
    .Y(_14179_));
 sky130_fd_sc_hd__o21ai_2 _24336_ (.A1(_13688_),
    .A2(_13690_),
    .B1(_14179_),
    .Y(_14180_));
 sky130_fd_sc_hd__or3_2 _24337_ (.A(_13688_),
    .B(_13690_),
    .C(_14179_),
    .X(_14181_));
 sky130_fd_sc_hd__o211ai_2 _24338_ (.A1(_14136_),
    .A2(_13740_),
    .B1(_14180_),
    .C1(_14181_),
    .Y(_14182_));
 sky130_fd_sc_hd__a211o_2 _24339_ (.A1(_14180_),
    .A2(_14181_),
    .B1(_14136_),
    .C1(_13740_),
    .X(_14183_));
 sky130_fd_sc_hd__nand4_2 _24340_ (.A(_14134_),
    .B(_14135_),
    .C(_14182_),
    .D(_14183_),
    .Y(_14184_));
 sky130_fd_sc_hd__a22o_2 _24341_ (.A1(_14134_),
    .A2(_14135_),
    .B1(_14182_),
    .B2(_14183_),
    .X(_14185_));
 sky130_fd_sc_hd__nand2_2 _24342_ (.A(_13696_),
    .B(_13747_),
    .Y(_14186_));
 sky130_fd_sc_hd__and3_2 _24343_ (.A(_14184_),
    .B(_14185_),
    .C(_14186_),
    .X(_14188_));
 sky130_fd_sc_hd__a21oi_2 _24344_ (.A1(_14184_),
    .A2(_14185_),
    .B1(_14186_),
    .Y(_14189_));
 sky130_fd_sc_hd__a211oi_2 _24345_ (.A1(_13743_),
    .A2(_13745_),
    .B1(_14188_),
    .C1(_14189_),
    .Y(_14190_));
 sky130_fd_sc_hd__o211a_2 _24346_ (.A1(_14188_),
    .A2(_14189_),
    .B1(_13743_),
    .C1(_13745_),
    .X(_14191_));
 sky130_fd_sc_hd__nor2_2 _24347_ (.A(_14190_),
    .B(_14191_),
    .Y(_14192_));
 sky130_fd_sc_hd__o21a_2 _24348_ (.A1(_13751_),
    .A2(_13753_),
    .B1(_14192_),
    .X(_14193_));
 sky130_fd_sc_hd__nor3_2 _24349_ (.A(_13751_),
    .B(_13753_),
    .C(_14192_),
    .Y(_14194_));
 sky130_fd_sc_hd__a211oi_2 _24350_ (.A1(_13711_),
    .A2(_13717_),
    .B1(_14193_),
    .C1(_14194_),
    .Y(_14195_));
 sky130_fd_sc_hd__o211a_2 _24351_ (.A1(_14193_),
    .A2(_14194_),
    .B1(_13711_),
    .C1(_13717_),
    .X(_14196_));
 sky130_fd_sc_hd__o211a_2 _24352_ (.A1(_14195_),
    .A2(_14196_),
    .B1(_13756_),
    .C1(_13759_),
    .X(_14197_));
 sky130_fd_sc_hd__a211o_2 _24353_ (.A1(_13756_),
    .A2(_13759_),
    .B1(_14195_),
    .C1(_14196_),
    .X(_14199_));
 sky130_fd_sc_hd__or2b_2 _24354_ (.A(_14197_),
    .B_N(_14199_),
    .X(_14200_));
 sky130_fd_sc_hd__inv_2 _24355_ (.A(_14200_),
    .Y(_14201_));
 sky130_fd_sc_hd__nand2_2 _24356_ (.A(_13765_),
    .B(_13767_),
    .Y(_14202_));
 sky130_fd_sc_hd__nand2_2 _24357_ (.A(_13763_),
    .B(_14202_),
    .Y(_14203_));
 sky130_fd_sc_hd__xnor2_2 _24358_ (.A(_14201_),
    .B(_14203_),
    .Y(_14204_));
 sky130_fd_sc_hd__o21ai_2 _24359_ (.A1(_14081_),
    .A2(_14082_),
    .B1(_14204_),
    .Y(_14205_));
 sky130_fd_sc_hd__or3_2 _24360_ (.A(_14081_),
    .B(_14082_),
    .C(_14204_),
    .X(_14206_));
 sky130_fd_sc_hd__nand2_2 _24361_ (.A(_14205_),
    .B(_14206_),
    .Y(_14207_));
 sky130_fd_sc_hd__a21o_2 _24362_ (.A1(_13640_),
    .A2(_13922_),
    .B1(_13921_),
    .X(_14208_));
 sky130_fd_sc_hd__xnor2_2 _24363_ (.A(_14207_),
    .B(_14208_),
    .Y(oO[43]));
 sky130_fd_sc_hd__inv_2 _24364_ (.A(_14206_),
    .Y(_14210_));
 sky130_fd_sc_hd__a211o_2 _24365_ (.A1(_13921_),
    .A2(_14205_),
    .B1(_14210_),
    .C1(_13638_),
    .X(_14211_));
 sky130_fd_sc_hd__nand2_2 _24366_ (.A(_13920_),
    .B(_14206_),
    .Y(_14212_));
 sky130_fd_sc_hd__a22oi_2 _24367_ (.A1(iY[14]),
    .A2(iX[30]),
    .B1(iX[31]),
    .B2(iY[13]),
    .Y(_14213_));
 sky130_fd_sc_hd__and3_2 _24368_ (.A(iY[14]),
    .B(iX[31]),
    .C(_13643_),
    .X(_14214_));
 sky130_fd_sc_hd__a21o_2 _24369_ (.A1(_14111_),
    .A2(_13680_),
    .B1(_14122_),
    .X(_14215_));
 sky130_fd_sc_hd__and4_2 _24370_ (.A(iY[21]),
    .B(iX[22]),
    .C(iY[22]),
    .D(iX[23]),
    .X(_14216_));
 sky130_fd_sc_hd__a22oi_2 _24371_ (.A1(iX[22]),
    .A2(iY[22]),
    .B1(iX[23]),
    .B2(iY[21]),
    .Y(_14217_));
 sky130_fd_sc_hd__nor2_2 _24372_ (.A(_14216_),
    .B(_14217_),
    .Y(_14218_));
 sky130_fd_sc_hd__nand2_2 _24373_ (.A(iX[21]),
    .B(iY[23]),
    .Y(_14220_));
 sky130_fd_sc_hd__xnor2_2 _24374_ (.A(_14218_),
    .B(_14220_),
    .Y(_14221_));
 sky130_fd_sc_hd__and4_2 _24375_ (.A(iY[18]),
    .B(iY[19]),
    .C(iX[25]),
    .D(iX[26]),
    .X(_14222_));
 sky130_fd_sc_hd__a22oi_2 _24376_ (.A1(iY[19]),
    .A2(iX[25]),
    .B1(iX[26]),
    .B2(iY[18]),
    .Y(_14223_));
 sky130_fd_sc_hd__nor2_2 _24377_ (.A(_14222_),
    .B(_14223_),
    .Y(_14224_));
 sky130_fd_sc_hd__nand2_2 _24378_ (.A(iY[20]),
    .B(iX[24]),
    .Y(_14225_));
 sky130_fd_sc_hd__xnor2_2 _24379_ (.A(_14224_),
    .B(_14225_),
    .Y(_14226_));
 sky130_fd_sc_hd__o21ba_2 _24380_ (.A1(_14101_),
    .A2(_14103_),
    .B1_N(_14100_),
    .X(_14227_));
 sky130_fd_sc_hd__xnor2_2 _24381_ (.A(_14226_),
    .B(_14227_),
    .Y(_14228_));
 sky130_fd_sc_hd__and2_2 _24382_ (.A(_14221_),
    .B(_14228_),
    .X(_14229_));
 sky130_fd_sc_hd__nor2_2 _24383_ (.A(_14221_),
    .B(_14228_),
    .Y(_14231_));
 sky130_fd_sc_hd__or2_2 _24384_ (.A(_14229_),
    .B(_14231_),
    .X(_14232_));
 sky130_fd_sc_hd__nand2_2 _24385_ (.A(_14112_),
    .B(_14120_),
    .Y(_14233_));
 sky130_fd_sc_hd__a31o_2 _24386_ (.A1(iY[17]),
    .A2(iX[26]),
    .A3(_14115_),
    .B1(_14113_),
    .X(_14234_));
 sky130_fd_sc_hd__and4_2 _24387_ (.A(iY[15]),
    .B(iY[16]),
    .C(iX[28]),
    .D(iX[29]),
    .X(_14235_));
 sky130_fd_sc_hd__a22oi_2 _24388_ (.A1(iY[16]),
    .A2(iX[28]),
    .B1(iX[29]),
    .B2(iY[15]),
    .Y(_14236_));
 sky130_fd_sc_hd__nor2_2 _24389_ (.A(_14235_),
    .B(_14236_),
    .Y(_14237_));
 sky130_fd_sc_hd__nand2_2 _24390_ (.A(iY[17]),
    .B(iX[27]),
    .Y(_14238_));
 sky130_fd_sc_hd__xnor2_2 _24391_ (.A(_14237_),
    .B(_14238_),
    .Y(_14239_));
 sky130_fd_sc_hd__o21ai_2 _24392_ (.A1(_14084_),
    .A2(_14086_),
    .B1(_14239_),
    .Y(_14240_));
 sky130_fd_sc_hd__or3_2 _24393_ (.A(_14084_),
    .B(_14086_),
    .C(_14239_),
    .X(_14242_));
 sky130_fd_sc_hd__and2_2 _24394_ (.A(_14240_),
    .B(_14242_),
    .X(_14243_));
 sky130_fd_sc_hd__xnor2_2 _24395_ (.A(_14234_),
    .B(_14243_),
    .Y(_14244_));
 sky130_fd_sc_hd__a21oi_2 _24396_ (.A1(_14118_),
    .A2(_14233_),
    .B1(_14244_),
    .Y(_14245_));
 sky130_fd_sc_hd__and3_2 _24397_ (.A(_14118_),
    .B(_14233_),
    .C(_14244_),
    .X(_14246_));
 sky130_fd_sc_hd__or3_2 _24398_ (.A(_14232_),
    .B(_14245_),
    .C(_14246_),
    .X(_14247_));
 sky130_fd_sc_hd__o21ai_2 _24399_ (.A1(_14245_),
    .A2(_14246_),
    .B1(_14232_),
    .Y(_14248_));
 sky130_fd_sc_hd__and3_2 _24400_ (.A(_14090_),
    .B(_14247_),
    .C(_14248_),
    .X(_14249_));
 sky130_fd_sc_hd__a21oi_2 _24401_ (.A1(_14247_),
    .A2(_14248_),
    .B1(_14090_),
    .Y(_14250_));
 sky130_fd_sc_hd__a211oi_2 _24402_ (.A1(_14215_),
    .A2(_14125_),
    .B1(_14249_),
    .C1(_14250_),
    .Y(_14251_));
 sky130_fd_sc_hd__o211a_2 _24403_ (.A1(_14249_),
    .A2(_14250_),
    .B1(_14215_),
    .C1(_14125_),
    .X(_14253_));
 sky130_fd_sc_hd__or4_2 _24404_ (.A(_14213_),
    .B(_14214_),
    .C(_14251_),
    .D(_14253_),
    .X(_14254_));
 sky130_fd_sc_hd__o22ai_2 _24405_ (.A1(_14213_),
    .A2(_14214_),
    .B1(_14251_),
    .B2(_14253_),
    .Y(_14255_));
 sky130_fd_sc_hd__nand3_2 _24406_ (.A(_14131_),
    .B(_14254_),
    .C(_14255_),
    .Y(_14256_));
 sky130_fd_sc_hd__a21o_2 _24407_ (.A1(_14254_),
    .A2(_14255_),
    .B1(_14131_),
    .X(_14257_));
 sky130_fd_sc_hd__inv_2 _24408_ (.A(_14177_),
    .Y(_14258_));
 sky130_fd_sc_hd__or2b_2 _24409_ (.A(_14127_),
    .B_N(_14129_),
    .X(_14259_));
 sky130_fd_sc_hd__inv_2 _24410_ (.A(_14259_),
    .Y(_14260_));
 sky130_fd_sc_hd__or2b_2 _24411_ (.A(_14144_),
    .B_N(_14142_),
    .X(_14261_));
 sky130_fd_sc_hd__and4_2 _24412_ (.A(iX[16]),
    .B(iX[17]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_14262_));
 sky130_fd_sc_hd__a22oi_2 _24413_ (.A1(iX[17]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[16]),
    .Y(_14264_));
 sky130_fd_sc_hd__nor2_2 _24414_ (.A(_14262_),
    .B(_14264_),
    .Y(_14265_));
 sky130_fd_sc_hd__nand2_2 _24415_ (.A(iX[15]),
    .B(iY[29]),
    .Y(_14266_));
 sky130_fd_sc_hd__xnor2_2 _24416_ (.A(_14265_),
    .B(_14266_),
    .Y(_14267_));
 sky130_fd_sc_hd__o21ba_2 _24417_ (.A1(_14139_),
    .A2(_14141_),
    .B1_N(_14138_),
    .X(_14268_));
 sky130_fd_sc_hd__xnor2_2 _24418_ (.A(_14267_),
    .B(_14268_),
    .Y(_14269_));
 sky130_fd_sc_hd__nand3_2 _24419_ (.A(iX[14]),
    .B(iY[30]),
    .C(_14269_),
    .Y(_14270_));
 sky130_fd_sc_hd__a21o_2 _24420_ (.A1(iX[14]),
    .A2(iY[30]),
    .B1(_14269_),
    .X(_14271_));
 sky130_fd_sc_hd__nand2_2 _24421_ (.A(_14270_),
    .B(_14271_),
    .Y(_14272_));
 sky130_fd_sc_hd__a21o_2 _24422_ (.A1(_14261_),
    .A2(_14146_),
    .B1(_14272_),
    .X(_14273_));
 sky130_fd_sc_hd__nand3_2 _24423_ (.A(_14261_),
    .B(_14146_),
    .C(_14272_),
    .Y(_14275_));
 sky130_fd_sc_hd__nand2_2 _24424_ (.A(_14273_),
    .B(_14275_),
    .Y(_14276_));
 sky130_fd_sc_hd__nand2_2 _24425_ (.A(iX[13]),
    .B(iY[31]),
    .Y(_14277_));
 sky130_fd_sc_hd__nand2_2 _24426_ (.A(_14276_),
    .B(_14277_),
    .Y(_14278_));
 sky130_fd_sc_hd__or2_2 _24427_ (.A(_14276_),
    .B(_14277_),
    .X(_14279_));
 sky130_fd_sc_hd__and2_2 _24428_ (.A(_14278_),
    .B(_14279_),
    .X(_14280_));
 sky130_fd_sc_hd__or2b_2 _24429_ (.A(_14160_),
    .B_N(_14166_),
    .X(_14281_));
 sky130_fd_sc_hd__or2b_2 _24430_ (.A(_14159_),
    .B_N(_14167_),
    .X(_14282_));
 sky130_fd_sc_hd__and2b_2 _24431_ (.A_N(_14105_),
    .B(_14104_),
    .X(_14283_));
 sky130_fd_sc_hd__o21ba_2 _24432_ (.A1(_14162_),
    .A2(_14164_),
    .B1_N(_14161_),
    .X(_14284_));
 sky130_fd_sc_hd__o21ba_2 _24433_ (.A1(_14095_),
    .A2(_14097_),
    .B1_N(_14094_),
    .X(_14286_));
 sky130_fd_sc_hd__and4_2 _24434_ (.A(iX[19]),
    .B(iX[20]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_14287_));
 sky130_fd_sc_hd__a22oi_2 _24435_ (.A1(iX[20]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[19]),
    .Y(_14288_));
 sky130_fd_sc_hd__nor2_2 _24436_ (.A(_14287_),
    .B(_14288_),
    .Y(_14289_));
 sky130_fd_sc_hd__nand2_2 _24437_ (.A(iX[18]),
    .B(iY[26]),
    .Y(_14290_));
 sky130_fd_sc_hd__xnor2_2 _24438_ (.A(_14289_),
    .B(_14290_),
    .Y(_14291_));
 sky130_fd_sc_hd__xnor2_2 _24439_ (.A(_14286_),
    .B(_14291_),
    .Y(_14292_));
 sky130_fd_sc_hd__xnor2_2 _24440_ (.A(_14284_),
    .B(_14292_),
    .Y(_14293_));
 sky130_fd_sc_hd__o21a_2 _24441_ (.A1(_14283_),
    .A2(_14107_),
    .B1(_14293_),
    .X(_14294_));
 sky130_fd_sc_hd__nor3_2 _24442_ (.A(_14283_),
    .B(_14107_),
    .C(_14293_),
    .Y(_14295_));
 sky130_fd_sc_hd__a211oi_2 _24443_ (.A1(_14281_),
    .A2(_14282_),
    .B1(_14294_),
    .C1(_14295_),
    .Y(_14297_));
 sky130_fd_sc_hd__o211a_2 _24444_ (.A1(_14294_),
    .A2(_14295_),
    .B1(_14281_),
    .C1(_14282_),
    .X(_14298_));
 sky130_fd_sc_hd__nor2_2 _24445_ (.A(_14169_),
    .B(_14171_),
    .Y(_14299_));
 sky130_fd_sc_hd__or3_2 _24446_ (.A(_14297_),
    .B(_14298_),
    .C(_14299_),
    .X(_14300_));
 sky130_fd_sc_hd__o21ai_2 _24447_ (.A1(_14297_),
    .A2(_14298_),
    .B1(_14299_),
    .Y(_14301_));
 sky130_fd_sc_hd__and3_2 _24448_ (.A(_14280_),
    .B(_14300_),
    .C(_14301_),
    .X(_14302_));
 sky130_fd_sc_hd__a21oi_2 _24449_ (.A1(_14300_),
    .A2(_14301_),
    .B1(_14280_),
    .Y(_14303_));
 sky130_fd_sc_hd__or3_2 _24450_ (.A(_14260_),
    .B(_14302_),
    .C(_14303_),
    .X(_14304_));
 sky130_fd_sc_hd__o21ai_2 _24451_ (.A1(_14302_),
    .A2(_14303_),
    .B1(_14260_),
    .Y(_14305_));
 sky130_fd_sc_hd__nand2_2 _24452_ (.A(_14304_),
    .B(_14305_),
    .Y(_14306_));
 sky130_fd_sc_hd__a21o_2 _24453_ (.A1(_14174_),
    .A2(_14258_),
    .B1(_14306_),
    .X(_14308_));
 sky130_fd_sc_hd__nand3_2 _24454_ (.A(_14174_),
    .B(_14258_),
    .C(_14306_),
    .Y(_14309_));
 sky130_fd_sc_hd__nand4_2 _24455_ (.A(_14256_),
    .B(_14257_),
    .C(_14308_),
    .D(_14309_),
    .Y(_14310_));
 sky130_fd_sc_hd__a22o_2 _24456_ (.A1(_14256_),
    .A2(_14257_),
    .B1(_14308_),
    .B2(_14309_),
    .X(_14311_));
 sky130_fd_sc_hd__nand2_2 _24457_ (.A(_14134_),
    .B(_14184_),
    .Y(_14312_));
 sky130_fd_sc_hd__and3_2 _24458_ (.A(_14310_),
    .B(_14311_),
    .C(_14312_),
    .X(_14313_));
 sky130_fd_sc_hd__a21oi_2 _24459_ (.A1(_14310_),
    .A2(_14311_),
    .B1(_14312_),
    .Y(_14314_));
 sky130_fd_sc_hd__or2_2 _24460_ (.A(_14313_),
    .B(_14314_),
    .X(_14315_));
 sky130_fd_sc_hd__nand2_2 _24461_ (.A(_14180_),
    .B(_14182_),
    .Y(_14316_));
 sky130_fd_sc_hd__xnor2_2 _24462_ (.A(_14315_),
    .B(_14316_),
    .Y(_14317_));
 sky130_fd_sc_hd__o21ai_2 _24463_ (.A1(_14188_),
    .A2(_14190_),
    .B1(_14317_),
    .Y(_14319_));
 sky130_fd_sc_hd__or3_2 _24464_ (.A(_14188_),
    .B(_14190_),
    .C(_14317_),
    .X(_14320_));
 sky130_fd_sc_hd__and2_2 _24465_ (.A(_14319_),
    .B(_14320_),
    .X(_14321_));
 sky130_fd_sc_hd__o21ai_2 _24466_ (.A1(_14149_),
    .A2(_14153_),
    .B1(_14321_),
    .Y(_14322_));
 sky130_fd_sc_hd__or3_2 _24467_ (.A(_14149_),
    .B(_14153_),
    .C(_14321_),
    .X(_14323_));
 sky130_fd_sc_hd__nand2_2 _24468_ (.A(_14322_),
    .B(_14323_),
    .Y(_14324_));
 sky130_fd_sc_hd__nor2_2 _24469_ (.A(_14193_),
    .B(_14195_),
    .Y(_14325_));
 sky130_fd_sc_hd__nor2_2 _24470_ (.A(_14324_),
    .B(_14325_),
    .Y(_14326_));
 sky130_fd_sc_hd__and2_2 _24471_ (.A(_14324_),
    .B(_14325_),
    .X(_14327_));
 sky130_fd_sc_hd__or2_2 _24472_ (.A(_14326_),
    .B(_14327_),
    .X(_14328_));
 sky130_fd_sc_hd__a311oi_2 _24473_ (.A1(_13763_),
    .A2(_14202_),
    .A3(_14199_),
    .B1(_14328_),
    .C1(_14197_),
    .Y(_14330_));
 sky130_fd_sc_hd__nand2_2 _24474_ (.A(_13765_),
    .B(_14201_),
    .Y(_14331_));
 sky130_fd_sc_hd__o221a_2 _24475_ (.A1(_13763_),
    .A2(_14197_),
    .B1(_14331_),
    .B2(_13766_),
    .C1(_14199_),
    .X(_14332_));
 sky130_fd_sc_hd__o311a_2 _24476_ (.A1(_13485_),
    .A2(_13483_),
    .A3(_14331_),
    .B1(_14332_),
    .C1(_14328_),
    .X(_14333_));
 sky130_fd_sc_hd__or2_2 _24477_ (.A(_14330_),
    .B(_14333_),
    .X(_14334_));
 sky130_fd_sc_hd__buf_1 _24478_ (.A(_14334_),
    .X(_14335_));
 sky130_fd_sc_hd__or3b_2 _24479_ (.A(_13984_),
    .B(_13985_),
    .C_N(_13986_),
    .X(_14336_));
 sky130_fd_sc_hd__o21bai_2 _24480_ (.A1(_13984_),
    .A2(_13985_),
    .B1_N(_13986_),
    .Y(_14337_));
 sky130_fd_sc_hd__nand4_2 _24481_ (.A(_13554_),
    .B(_13906_),
    .C(_14336_),
    .D(_14337_),
    .Y(_14338_));
 sky130_fd_sc_hd__and3_2 _24482_ (.A(_13904_),
    .B(_14336_),
    .C(_14337_),
    .X(_14339_));
 sky130_fd_sc_hd__a2bb2o_2 _24483_ (.A1_N(_13954_),
    .A2_N(_13956_),
    .B1(_13866_),
    .B2(_13953_),
    .X(_14341_));
 sky130_fd_sc_hd__o21ai_2 _24484_ (.A1(_13929_),
    .A2(_13930_),
    .B1(_13927_),
    .Y(_14342_));
 sky130_fd_sc_hd__buf_1 _24485_ (.A(_13231_),
    .X(_14343_));
 sky130_fd_sc_hd__nor2_2 _24486_ (.A(_14343_),
    .B(_12772_),
    .Y(_14344_));
 sky130_fd_sc_hd__xnor2_2 _24487_ (.A(_13953_),
    .B(_14344_),
    .Y(_14345_));
 sky130_fd_sc_hd__buf_6 _24488_ (.A(_12223_),
    .X(_14346_));
 sky130_fd_sc_hd__nor2_2 _24489_ (.A(_14346_),
    .B(_13273_),
    .Y(_14347_));
 sky130_fd_sc_hd__xnor2_2 _24490_ (.A(_14345_),
    .B(_14347_),
    .Y(_14348_));
 sky130_fd_sc_hd__xnor2_2 _24491_ (.A(_14342_),
    .B(_14348_),
    .Y(_14349_));
 sky130_fd_sc_hd__xnor2_2 _24492_ (.A(_14341_),
    .B(_14349_),
    .Y(_14350_));
 sky130_fd_sc_hd__buf_1 _24493_ (.A(_13241_),
    .X(_14352_));
 sky130_fd_sc_hd__or4_2 _24494_ (.A(_13926_),
    .B(_12248_),
    .C(_14352_),
    .D(_13502_),
    .X(_14353_));
 sky130_fd_sc_hd__a22o_2 _24495_ (.A1(_12242_),
    .A2(_13244_),
    .B1(_13496_),
    .B2(_11842_),
    .X(_14354_));
 sky130_fd_sc_hd__nand2_2 _24496_ (.A(_14353_),
    .B(_14354_),
    .Y(_14355_));
 sky130_fd_sc_hd__xnor2_2 _24497_ (.A(_12474_),
    .B(_12476_),
    .Y(_14356_));
 sky130_fd_sc_hd__buf_1 _24498_ (.A(_12808_),
    .X(_14357_));
 sky130_fd_sc_hd__nor2_2 _24499_ (.A(_14356_),
    .B(_14357_),
    .Y(_14358_));
 sky130_fd_sc_hd__xnor2_2 _24500_ (.A(_14355_),
    .B(_14358_),
    .Y(_14359_));
 sky130_fd_sc_hd__nor2_2 _24501_ (.A(_11793_),
    .B(_13842_),
    .Y(_14360_));
 sky130_fd_sc_hd__nor2_2 _24502_ (.A(_11566_),
    .B(_13934_),
    .Y(_14361_));
 sky130_fd_sc_hd__nor2_2 _24503_ (.A(iX[11]),
    .B(iX[43]),
    .Y(_14363_));
 sky130_fd_sc_hd__xnor2_2 _24504_ (.A(iX[12]),
    .B(iX[44]),
    .Y(_14364_));
 sky130_fd_sc_hd__a21o_2 _24505_ (.A1(iX[11]),
    .A2(iX[43]),
    .B1(_13835_),
    .X(_14365_));
 sky130_fd_sc_hd__a21oi_2 _24506_ (.A1(_13838_),
    .A2(_13841_),
    .B1(_14365_),
    .Y(_14366_));
 sky130_fd_sc_hd__or3_2 _24507_ (.A(_14363_),
    .B(_14364_),
    .C(_14366_),
    .X(_14367_));
 sky130_fd_sc_hd__o21ai_2 _24508_ (.A1(_14363_),
    .A2(_14366_),
    .B1(_14364_),
    .Y(_14368_));
 sky130_fd_sc_hd__and3_2 _24509_ (.A(_11583_),
    .B(_14367_),
    .C(_14368_),
    .X(_14369_));
 sky130_fd_sc_hd__a32o_2 _24510_ (.A1(_11379_),
    .A2(_14367_),
    .A3(_14368_),
    .B1(_11583_),
    .B2(_13937_),
    .X(_14370_));
 sky130_fd_sc_hd__a21boi_2 _24511_ (.A1(_14361_),
    .A2(_14369_),
    .B1_N(_14370_),
    .Y(_14371_));
 sky130_fd_sc_hd__xnor2_2 _24512_ (.A(_14360_),
    .B(_14371_),
    .Y(_14372_));
 sky130_fd_sc_hd__and2_2 _24513_ (.A(_13936_),
    .B(_13940_),
    .X(_14374_));
 sky130_fd_sc_hd__xor2_2 _24514_ (.A(_14372_),
    .B(_14374_),
    .X(_14375_));
 sky130_fd_sc_hd__xnor2_2 _24515_ (.A(_14359_),
    .B(_14375_),
    .Y(_14376_));
 sky130_fd_sc_hd__and2_2 _24516_ (.A(_13943_),
    .B(_13945_),
    .X(_14377_));
 sky130_fd_sc_hd__xor2_2 _24517_ (.A(_14376_),
    .B(_14377_),
    .X(_14378_));
 sky130_fd_sc_hd__xnor2_2 _24518_ (.A(_14350_),
    .B(_14378_),
    .Y(_14379_));
 sky130_fd_sc_hd__and2_2 _24519_ (.A(_13949_),
    .B(_13961_),
    .X(_14380_));
 sky130_fd_sc_hd__xor2_2 _24520_ (.A(_14379_),
    .B(_14380_),
    .X(_14381_));
 sky130_fd_sc_hd__or2_2 _24521_ (.A(_13894_),
    .B(_13974_),
    .X(_14382_));
 sky130_fd_sc_hd__and2b_2 _24522_ (.A_N(_13959_),
    .B(_13951_),
    .X(_14383_));
 sky130_fd_sc_hd__a21o_2 _24523_ (.A1(_13952_),
    .A2(_13958_),
    .B1(_14383_),
    .X(_14385_));
 sky130_fd_sc_hd__xnor2_2 _24524_ (.A(_13538_),
    .B(_13540_),
    .Y(_14386_));
 sky130_fd_sc_hd__or4_2 _24525_ (.A(_12468_),
    .B(_11827_),
    .C(_14386_),
    .D(_13891_),
    .X(_14387_));
 sky130_fd_sc_hd__buf_1 _24526_ (.A(_11829_),
    .X(_14388_));
 sky130_fd_sc_hd__a22o_2 _24527_ (.A1(_14388_),
    .A2(_13543_),
    .B1(_13888_),
    .B2(_12827_),
    .X(_14389_));
 sky130_fd_sc_hd__nand2_2 _24528_ (.A(_14387_),
    .B(_14389_),
    .Y(_14390_));
 sky130_fd_sc_hd__xnor2_2 _24529_ (.A(_13970_),
    .B(_13971_),
    .Y(_14391_));
 sky130_fd_sc_hd__buf_1 _24530_ (.A(_14391_),
    .X(_14392_));
 sky130_fd_sc_hd__nand2_2 _24531_ (.A(_12838_),
    .B(_14392_),
    .Y(_14393_));
 sky130_fd_sc_hd__xnor2_2 _24532_ (.A(_14390_),
    .B(_14393_),
    .Y(_14394_));
 sky130_fd_sc_hd__a21oi_2 _24533_ (.A1(_13968_),
    .A2(_13973_),
    .B1(_13967_),
    .Y(_14396_));
 sky130_fd_sc_hd__xor2_2 _24534_ (.A(_14394_),
    .B(_14396_),
    .X(_14397_));
 sky130_fd_sc_hd__nor4bb_2 _24535_ (.A(_13884_),
    .B(_13970_),
    .C_N(_13885_),
    .D_N(_13536_),
    .Y(_14398_));
 sky130_fd_sc_hd__o211a_2 _24536_ (.A1(iY[11]),
    .A2(iY[43]),
    .B1(iY[42]),
    .C1(iY[10]),
    .X(_14399_));
 sky130_fd_sc_hd__a211o_2 _24537_ (.A1(iY[11]),
    .A2(iY[43]),
    .B1(_14398_),
    .C1(_14399_),
    .X(_14400_));
 sky130_fd_sc_hd__and4bb_2 _24538_ (.A_N(_13884_),
    .B_N(_13970_),
    .C(_13536_),
    .D(_13537_),
    .X(_14401_));
 sky130_fd_sc_hd__o2111a_2 _24539_ (.A1(_12771_),
    .A2(_13269_),
    .B1(_13271_),
    .C1(_14401_),
    .D1(_13267_),
    .X(_14402_));
 sky130_fd_sc_hd__nand2_2 _24540_ (.A(iY[12]),
    .B(iY[44]),
    .Y(_14403_));
 sky130_fd_sc_hd__or2_2 _24541_ (.A(iY[12]),
    .B(iY[44]),
    .X(_14404_));
 sky130_fd_sc_hd__nand2_2 _24542_ (.A(_14403_),
    .B(_14404_),
    .Y(_14405_));
 sky130_fd_sc_hd__o21bai_2 _24543_ (.A1(_14400_),
    .A2(_14402_),
    .B1_N(_14405_),
    .Y(_14407_));
 sky130_fd_sc_hd__or3b_2 _24544_ (.A(_14400_),
    .B(_14402_),
    .C_N(_14405_),
    .X(_14408_));
 sky130_fd_sc_hd__and2_2 _24545_ (.A(_14407_),
    .B(_14408_),
    .X(_14409_));
 sky130_fd_sc_hd__buf_1 _24546_ (.A(_14409_),
    .X(_14410_));
 sky130_fd_sc_hd__buf_1 _24547_ (.A(_14410_),
    .X(_14411_));
 sky130_fd_sc_hd__nand2_2 _24548_ (.A(_11374_),
    .B(_14411_),
    .Y(_14412_));
 sky130_fd_sc_hd__xnor2_2 _24549_ (.A(_14397_),
    .B(_14412_),
    .Y(_14413_));
 sky130_fd_sc_hd__xnor2_2 _24550_ (.A(_14385_),
    .B(_14413_),
    .Y(_14414_));
 sky130_fd_sc_hd__xor2_2 _24551_ (.A(_14382_),
    .B(_14414_),
    .X(_14415_));
 sky130_fd_sc_hd__xor2_2 _24552_ (.A(_14381_),
    .B(_14415_),
    .X(_14416_));
 sky130_fd_sc_hd__nor2_2 _24553_ (.A(_13964_),
    .B(_13980_),
    .Y(_14418_));
 sky130_fd_sc_hd__xnor2_2 _24554_ (.A(_14416_),
    .B(_14418_),
    .Y(_14419_));
 sky130_fd_sc_hd__xnor2_2 _24555_ (.A(_13976_),
    .B(_14419_),
    .Y(_14420_));
 sky130_fd_sc_hd__a21boi_2 _24556_ (.A1(_13923_),
    .A2(_13983_),
    .B1_N(_13982_),
    .Y(_14421_));
 sky130_fd_sc_hd__xnor2_2 _24557_ (.A(_14420_),
    .B(_14421_),
    .Y(_14422_));
 sky130_fd_sc_hd__xnor2_2 _24558_ (.A(_13987_),
    .B(_14422_),
    .Y(_14423_));
 sky130_fd_sc_hd__xnor2_2 _24559_ (.A(_14339_),
    .B(_14423_),
    .Y(_14424_));
 sky130_fd_sc_hd__xor2_2 _24560_ (.A(_14338_),
    .B(_14424_),
    .X(_14425_));
 sky130_fd_sc_hd__nand2b_2 _24561_ (.A_N(_13994_),
    .B(_13997_),
    .Y(_14426_));
 sky130_fd_sc_hd__xor2_2 _24562_ (.A(_14425_),
    .B(_14426_),
    .X(_14427_));
 sky130_fd_sc_hd__nor3_2 _24563_ (.A(_13822_),
    .B(_13821_),
    .C(_14060_),
    .Y(_14429_));
 sky130_fd_sc_hd__nand2_2 _24564_ (.A(_14056_),
    .B(_14059_),
    .Y(_14430_));
 sky130_fd_sc_hd__nand2_2 _24565_ (.A(_14004_),
    .B(_14005_),
    .Y(_14431_));
 sky130_fd_sc_hd__nand2_2 _24566_ (.A(_14006_),
    .B(_14012_),
    .Y(_14432_));
 sky130_fd_sc_hd__and4_2 _24567_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[41]),
    .D(iX[42]),
    .X(_14433_));
 sky130_fd_sc_hd__a22oi_2 _24568_ (.A1(iY[35]),
    .A2(iX[41]),
    .B1(iX[42]),
    .B2(iY[34]),
    .Y(_14434_));
 sky130_fd_sc_hd__nor2_2 _24569_ (.A(_14433_),
    .B(_14434_),
    .Y(_14435_));
 sky130_fd_sc_hd__nand2_2 _24570_ (.A(iY[33]),
    .B(iX[43]),
    .Y(_14436_));
 sky130_fd_sc_hd__xnor2_2 _24571_ (.A(_14435_),
    .B(_14436_),
    .Y(_14437_));
 sky130_fd_sc_hd__o21ba_2 _24572_ (.A1(_14001_),
    .A2(_14003_),
    .B1_N(_13999_),
    .X(_14438_));
 sky130_fd_sc_hd__xnor2_2 _24573_ (.A(_14437_),
    .B(_14438_),
    .Y(_14440_));
 sky130_fd_sc_hd__and4_2 _24574_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[40]),
    .D(iX[44]),
    .X(_14441_));
 sky130_fd_sc_hd__a22oi_2 _24575_ (.A1(iY[36]),
    .A2(iX[40]),
    .B1(iX[44]),
    .B2(iY[32]),
    .Y(_14442_));
 sky130_fd_sc_hd__nor2_2 _24576_ (.A(_14441_),
    .B(_14442_),
    .Y(_14443_));
 sky130_fd_sc_hd__nand2_2 _24577_ (.A(iY[37]),
    .B(iX[39]),
    .Y(_14444_));
 sky130_fd_sc_hd__xnor2_2 _24578_ (.A(_14443_),
    .B(_14444_),
    .Y(_14445_));
 sky130_fd_sc_hd__xnor2_2 _24579_ (.A(_14440_),
    .B(_14445_),
    .Y(_14446_));
 sky130_fd_sc_hd__a21o_2 _24580_ (.A1(_14431_),
    .A2(_14432_),
    .B1(_14446_),
    .X(_14447_));
 sky130_fd_sc_hd__nand3_2 _24581_ (.A(_14431_),
    .B(_14432_),
    .C(_14446_),
    .Y(_14448_));
 sky130_fd_sc_hd__o21ba_2 _24582_ (.A1(_14019_),
    .A2(_14021_),
    .B1_N(_14018_),
    .X(_14449_));
 sky130_fd_sc_hd__o21ba_2 _24583_ (.A1(_14008_),
    .A2(_14010_),
    .B1_N(_14007_),
    .X(_14451_));
 sky130_fd_sc_hd__and4_2 _24584_ (.A(iX[37]),
    .B(iX[38]),
    .C(iY[38]),
    .D(iY[39]),
    .X(_14452_));
 sky130_fd_sc_hd__a22oi_2 _24585_ (.A1(iX[38]),
    .A2(iY[38]),
    .B1(iY[39]),
    .B2(iX[37]),
    .Y(_14453_));
 sky130_fd_sc_hd__nor2_2 _24586_ (.A(_14452_),
    .B(_14453_),
    .Y(_14454_));
 sky130_fd_sc_hd__nand2_2 _24587_ (.A(iX[36]),
    .B(iY[40]),
    .Y(_14455_));
 sky130_fd_sc_hd__xnor2_2 _24588_ (.A(_14454_),
    .B(_14455_),
    .Y(_14456_));
 sky130_fd_sc_hd__xnor2_2 _24589_ (.A(_14451_),
    .B(_14456_),
    .Y(_14457_));
 sky130_fd_sc_hd__xnor2_2 _24590_ (.A(_14449_),
    .B(_14457_),
    .Y(_14458_));
 sky130_fd_sc_hd__and3_2 _24591_ (.A(_14447_),
    .B(_14448_),
    .C(_14458_),
    .X(_14459_));
 sky130_fd_sc_hd__a21oi_2 _24592_ (.A1(_14447_),
    .A2(_14448_),
    .B1(_14458_),
    .Y(_14460_));
 sky130_fd_sc_hd__or2_2 _24593_ (.A(_14459_),
    .B(_14460_),
    .X(_14462_));
 sky130_fd_sc_hd__a21oi_2 _24594_ (.A1(_14014_),
    .A2(_14028_),
    .B1(_14462_),
    .Y(_14463_));
 sky130_fd_sc_hd__and3_2 _24595_ (.A(_14014_),
    .B(_14028_),
    .C(_14462_),
    .X(_14464_));
 sky130_fd_sc_hd__or2b_2 _24596_ (.A(_14016_),
    .B_N(_14026_),
    .X(_14465_));
 sky130_fd_sc_hd__nand2_2 _24597_ (.A(_14024_),
    .B(_14465_),
    .Y(_14466_));
 sky130_fd_sc_hd__and4_2 _24598_ (.A(iX[34]),
    .B(iX[35]),
    .C(iY[41]),
    .D(iY[42]),
    .X(_14467_));
 sky130_fd_sc_hd__a22oi_2 _24599_ (.A1(iX[35]),
    .A2(iY[41]),
    .B1(iY[42]),
    .B2(iX[34]),
    .Y(_14468_));
 sky130_fd_sc_hd__nor2_2 _24600_ (.A(_14467_),
    .B(_14468_),
    .Y(_14469_));
 sky130_fd_sc_hd__nand2_2 _24601_ (.A(iX[33]),
    .B(iY[43]),
    .Y(_14470_));
 sky130_fd_sc_hd__xnor2_2 _24602_ (.A(_14469_),
    .B(_14470_),
    .Y(_14471_));
 sky130_fd_sc_hd__o21ba_2 _24603_ (.A1(_14037_),
    .A2(_14039_),
    .B1_N(_14036_),
    .X(_14473_));
 sky130_fd_sc_hd__xnor2_2 _24604_ (.A(_14471_),
    .B(_14473_),
    .Y(_14474_));
 sky130_fd_sc_hd__nand3_2 _24605_ (.A(iX[32]),
    .B(iY[44]),
    .C(_14474_),
    .Y(_14475_));
 sky130_fd_sc_hd__a21o_2 _24606_ (.A1(iX[32]),
    .A2(iY[44]),
    .B1(_14474_),
    .X(_14476_));
 sky130_fd_sc_hd__nand2_2 _24607_ (.A(_14475_),
    .B(_14476_),
    .Y(_14477_));
 sky130_fd_sc_hd__xnor2_2 _24608_ (.A(_14466_),
    .B(_14477_),
    .Y(_14478_));
 sky130_fd_sc_hd__xnor2_2 _24609_ (.A(_14041_),
    .B(_14478_),
    .Y(_14479_));
 sky130_fd_sc_hd__or3_2 _24610_ (.A(_14463_),
    .B(_14464_),
    .C(_14479_),
    .X(_14480_));
 sky130_fd_sc_hd__o21ai_2 _24611_ (.A1(_14463_),
    .A2(_14464_),
    .B1(_14479_),
    .Y(_14481_));
 sky130_fd_sc_hd__nand2_2 _24612_ (.A(_14031_),
    .B(_14048_),
    .Y(_14482_));
 sky130_fd_sc_hd__nand3_2 _24613_ (.A(_14480_),
    .B(_14481_),
    .C(_14482_),
    .Y(_14484_));
 sky130_fd_sc_hd__a21o_2 _24614_ (.A1(_14480_),
    .A2(_14481_),
    .B1(_14482_),
    .X(_14485_));
 sky130_fd_sc_hd__and3_2 _24615_ (.A(_14045_),
    .B(_14484_),
    .C(_14485_),
    .X(_14486_));
 sky130_fd_sc_hd__a21oi_2 _24616_ (.A1(_14484_),
    .A2(_14485_),
    .B1(_14045_),
    .Y(_14487_));
 sky130_fd_sc_hd__a211oi_2 _24617_ (.A1(_14051_),
    .A2(_14054_),
    .B1(_14486_),
    .C1(_14487_),
    .Y(_14488_));
 sky130_fd_sc_hd__o211a_2 _24618_ (.A1(_14486_),
    .A2(_14487_),
    .B1(_14051_),
    .C1(_14054_),
    .X(_14489_));
 sky130_fd_sc_hd__or3_2 _24619_ (.A(_14430_),
    .B(_14488_),
    .C(_14489_),
    .X(_14490_));
 sky130_fd_sc_hd__o21ai_2 _24620_ (.A1(_14488_),
    .A2(_14489_),
    .B1(_14430_),
    .Y(_14491_));
 sky130_fd_sc_hd__or4bb_2 _24621_ (.A(_14061_),
    .B(_14060_),
    .C_N(_14490_),
    .D_N(_14491_),
    .X(_14492_));
 sky130_fd_sc_hd__a2bb2o_2 _24622_ (.A1_N(_14061_),
    .A2_N(_14060_),
    .B1(_14490_),
    .B2(_14491_),
    .X(_14493_));
 sky130_fd_sc_hd__and3_2 _24623_ (.A(_14429_),
    .B(_14492_),
    .C(_14493_),
    .X(_14495_));
 sky130_fd_sc_hd__a21oi_2 _24624_ (.A1(_14492_),
    .A2(_14493_),
    .B1(_14429_),
    .Y(_14496_));
 sky130_fd_sc_hd__or2_2 _24625_ (.A(_14495_),
    .B(_14496_),
    .X(_14497_));
 sky130_fd_sc_hd__a21boi_2 _24626_ (.A1(_14065_),
    .A2(_14069_),
    .B1_N(_14064_),
    .Y(_14498_));
 sky130_fd_sc_hd__xnor2_2 _24627_ (.A(_14497_),
    .B(_14498_),
    .Y(_14499_));
 sky130_fd_sc_hd__xor2_2 _24628_ (.A(_14427_),
    .B(_14499_),
    .X(_14500_));
 sky130_fd_sc_hd__xor2_2 _24629_ (.A(oO[12]),
    .B(_14500_),
    .X(_14501_));
 sky130_fd_sc_hd__o21ba_2 _24630_ (.A1(oO[11]),
    .A2(_14072_),
    .B1_N(_14071_),
    .X(_14502_));
 sky130_fd_sc_hd__xor2_2 _24631_ (.A(_14501_),
    .B(_14502_),
    .X(_14503_));
 sky130_fd_sc_hd__or2b_2 _24632_ (.A(_14074_),
    .B_N(_14076_),
    .X(_14504_));
 sky130_fd_sc_hd__o21ai_2 _24633_ (.A1(_14078_),
    .A2(_14080_),
    .B1(_14504_),
    .Y(_14506_));
 sky130_fd_sc_hd__xor2_2 _24634_ (.A(_14503_),
    .B(_14506_),
    .X(_14507_));
 sky130_fd_sc_hd__xor2_2 _24635_ (.A(_14335_),
    .B(_14507_),
    .X(_14508_));
 sky130_fd_sc_hd__inv_2 _24636_ (.A(_14508_),
    .Y(_14509_));
 sky130_fd_sc_hd__o2111a_2 _24637_ (.A1(_13637_),
    .A2(_14211_),
    .B1(_14212_),
    .C1(_14509_),
    .D1(_14205_),
    .X(_14510_));
 sky130_fd_sc_hd__o211ai_2 _24638_ (.A1(_13637_),
    .A2(_14211_),
    .B1(_14212_),
    .C1(_14205_),
    .Y(_14511_));
 sky130_fd_sc_hd__and2_2 _24639_ (.A(_14508_),
    .B(_14511_),
    .X(_14512_));
 sky130_fd_sc_hd__nor2_2 _24640_ (.A(_14510_),
    .B(_14512_),
    .Y(oO[44]));
 sky130_fd_sc_hd__o21bai_2 _24641_ (.A1(_14496_),
    .A2(_14498_),
    .B1_N(_14495_),
    .Y(_14513_));
 sky130_fd_sc_hd__inv_2 _24642_ (.A(_14488_),
    .Y(_14514_));
 sky130_fd_sc_hd__nor3_2 _24643_ (.A(_14463_),
    .B(_14464_),
    .C(_14479_),
    .Y(_14516_));
 sky130_fd_sc_hd__or2b_2 _24644_ (.A(_14438_),
    .B_N(_14437_),
    .X(_14517_));
 sky130_fd_sc_hd__nand2_2 _24645_ (.A(_14440_),
    .B(_14445_),
    .Y(_14518_));
 sky130_fd_sc_hd__and4_2 _24646_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[42]),
    .D(iX[43]),
    .X(_14519_));
 sky130_fd_sc_hd__a22oi_2 _24647_ (.A1(iY[35]),
    .A2(iX[42]),
    .B1(iX[43]),
    .B2(iY[34]),
    .Y(_14520_));
 sky130_fd_sc_hd__nor2_2 _24648_ (.A(_14519_),
    .B(_14520_),
    .Y(_14521_));
 sky130_fd_sc_hd__nand2_2 _24649_ (.A(iY[33]),
    .B(iX[44]),
    .Y(_14522_));
 sky130_fd_sc_hd__xnor2_2 _24650_ (.A(_14521_),
    .B(_14522_),
    .Y(_14523_));
 sky130_fd_sc_hd__o21ba_2 _24651_ (.A1(_14434_),
    .A2(_14436_),
    .B1_N(_14433_),
    .X(_14524_));
 sky130_fd_sc_hd__xnor2_2 _24652_ (.A(_14523_),
    .B(_14524_),
    .Y(_14525_));
 sky130_fd_sc_hd__and4_2 _24653_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[41]),
    .D(iX[45]),
    .X(_14527_));
 sky130_fd_sc_hd__a22oi_2 _24654_ (.A1(iY[36]),
    .A2(iX[41]),
    .B1(iX[45]),
    .B2(iY[32]),
    .Y(_14528_));
 sky130_fd_sc_hd__nor2_2 _24655_ (.A(_14527_),
    .B(_14528_),
    .Y(_14529_));
 sky130_fd_sc_hd__nand2_2 _24656_ (.A(iY[37]),
    .B(iX[40]),
    .Y(_14530_));
 sky130_fd_sc_hd__xnor2_2 _24657_ (.A(_14529_),
    .B(_14530_),
    .Y(_14531_));
 sky130_fd_sc_hd__xnor2_2 _24658_ (.A(_14525_),
    .B(_14531_),
    .Y(_14532_));
 sky130_fd_sc_hd__a21o_2 _24659_ (.A1(_14517_),
    .A2(_14518_),
    .B1(_14532_),
    .X(_14533_));
 sky130_fd_sc_hd__nand3_2 _24660_ (.A(_14517_),
    .B(_14518_),
    .C(_14532_),
    .Y(_14534_));
 sky130_fd_sc_hd__o21ba_2 _24661_ (.A1(_14453_),
    .A2(_14455_),
    .B1_N(_14452_),
    .X(_14535_));
 sky130_fd_sc_hd__o21ba_2 _24662_ (.A1(_14442_),
    .A2(_14444_),
    .B1_N(_14441_),
    .X(_14536_));
 sky130_fd_sc_hd__and4_2 _24663_ (.A(iX[38]),
    .B(iY[38]),
    .C(iX[39]),
    .D(iY[39]),
    .X(_14538_));
 sky130_fd_sc_hd__a22oi_2 _24664_ (.A1(iY[38]),
    .A2(iX[39]),
    .B1(iY[39]),
    .B2(iX[38]),
    .Y(_14539_));
 sky130_fd_sc_hd__nor2_2 _24665_ (.A(_14538_),
    .B(_14539_),
    .Y(_14540_));
 sky130_fd_sc_hd__nand2_2 _24666_ (.A(iX[37]),
    .B(iY[40]),
    .Y(_14541_));
 sky130_fd_sc_hd__xnor2_2 _24667_ (.A(_14540_),
    .B(_14541_),
    .Y(_14542_));
 sky130_fd_sc_hd__xnor2_2 _24668_ (.A(_14536_),
    .B(_14542_),
    .Y(_14543_));
 sky130_fd_sc_hd__xnor2_2 _24669_ (.A(_14535_),
    .B(_14543_),
    .Y(_14544_));
 sky130_fd_sc_hd__nand3_2 _24670_ (.A(_14533_),
    .B(_14534_),
    .C(_14544_),
    .Y(_14545_));
 sky130_fd_sc_hd__a21o_2 _24671_ (.A1(_14533_),
    .A2(_14534_),
    .B1(_14544_),
    .X(_14546_));
 sky130_fd_sc_hd__and2_2 _24672_ (.A(_14545_),
    .B(_14546_),
    .X(_14547_));
 sky130_fd_sc_hd__a21bo_2 _24673_ (.A1(_14448_),
    .A2(_14458_),
    .B1_N(_14447_),
    .X(_14549_));
 sky130_fd_sc_hd__xnor2_2 _24674_ (.A(_14547_),
    .B(_14549_),
    .Y(_14550_));
 sky130_fd_sc_hd__or2b_2 _24675_ (.A(_14473_),
    .B_N(_14471_),
    .X(_14551_));
 sky130_fd_sc_hd__and2b_2 _24676_ (.A_N(_14451_),
    .B(_14456_),
    .X(_14552_));
 sky130_fd_sc_hd__and2b_2 _24677_ (.A_N(_14449_),
    .B(_14457_),
    .X(_14553_));
 sky130_fd_sc_hd__a22oi_2 _24678_ (.A1(iX[33]),
    .A2(iY[44]),
    .B1(iY[45]),
    .B2(iX[32]),
    .Y(_14554_));
 sky130_fd_sc_hd__and4_2 _24679_ (.A(iX[33]),
    .B(iX[32]),
    .C(iY[44]),
    .D(iY[45]),
    .X(_14555_));
 sky130_fd_sc_hd__or2_2 _24680_ (.A(_14554_),
    .B(_14555_),
    .X(_14556_));
 sky130_fd_sc_hd__and4_2 _24681_ (.A(iX[35]),
    .B(iX[36]),
    .C(iY[41]),
    .D(iY[42]),
    .X(_14557_));
 sky130_fd_sc_hd__a22oi_2 _24682_ (.A1(iX[36]),
    .A2(iY[41]),
    .B1(iY[42]),
    .B2(iX[35]),
    .Y(_14558_));
 sky130_fd_sc_hd__nor2_2 _24683_ (.A(_14557_),
    .B(_14558_),
    .Y(_14560_));
 sky130_fd_sc_hd__nand2_2 _24684_ (.A(iX[34]),
    .B(iY[43]),
    .Y(_14561_));
 sky130_fd_sc_hd__xnor2_2 _24685_ (.A(_14560_),
    .B(_14561_),
    .Y(_14562_));
 sky130_fd_sc_hd__o21ba_2 _24686_ (.A1(_14468_),
    .A2(_14470_),
    .B1_N(_14467_),
    .X(_14563_));
 sky130_fd_sc_hd__xnor2_2 _24687_ (.A(_14562_),
    .B(_14563_),
    .Y(_14564_));
 sky130_fd_sc_hd__xnor2_2 _24688_ (.A(_14556_),
    .B(_14564_),
    .Y(_14565_));
 sky130_fd_sc_hd__o21a_2 _24689_ (.A1(_14552_),
    .A2(_14553_),
    .B1(_14565_),
    .X(_14566_));
 sky130_fd_sc_hd__nor3_2 _24690_ (.A(_14552_),
    .B(_14553_),
    .C(_14565_),
    .Y(_14567_));
 sky130_fd_sc_hd__a211oi_2 _24691_ (.A1(_14551_),
    .A2(_14475_),
    .B1(_14566_),
    .C1(_14567_),
    .Y(_14568_));
 sky130_fd_sc_hd__o211a_2 _24692_ (.A1(_14566_),
    .A2(_14567_),
    .B1(_14551_),
    .C1(_14475_),
    .X(_14569_));
 sky130_fd_sc_hd__or3_2 _24693_ (.A(_14550_),
    .B(_14568_),
    .C(_14569_),
    .X(_14571_));
 sky130_fd_sc_hd__o21ai_2 _24694_ (.A1(_14568_),
    .A2(_14569_),
    .B1(_14550_),
    .Y(_14572_));
 sky130_fd_sc_hd__o211a_2 _24695_ (.A1(_14463_),
    .A2(_14516_),
    .B1(_14571_),
    .C1(_14572_),
    .X(_14573_));
 sky130_fd_sc_hd__a211oi_2 _24696_ (.A1(_14571_),
    .A2(_14572_),
    .B1(_14463_),
    .C1(_14516_),
    .Y(_14574_));
 sky130_fd_sc_hd__nor2_2 _24697_ (.A(_14573_),
    .B(_14574_),
    .Y(_14575_));
 sky130_fd_sc_hd__a32oi_2 _24698_ (.A1(_14466_),
    .A2(_14475_),
    .A3(_14476_),
    .B1(_14478_),
    .B2(_14041_),
    .Y(_14576_));
 sky130_fd_sc_hd__xnor2_2 _24699_ (.A(_14575_),
    .B(_14576_),
    .Y(_14577_));
 sky130_fd_sc_hd__inv_2 _24700_ (.A(_14484_),
    .Y(_14578_));
 sky130_fd_sc_hd__nor2_2 _24701_ (.A(_14578_),
    .B(_14486_),
    .Y(_14579_));
 sky130_fd_sc_hd__xor2_2 _24702_ (.A(_14577_),
    .B(_14579_),
    .X(_14580_));
 sky130_fd_sc_hd__or2_2 _24703_ (.A(_14514_),
    .B(_14580_),
    .X(_14581_));
 sky130_fd_sc_hd__nand2_2 _24704_ (.A(_14514_),
    .B(_14580_),
    .Y(_14582_));
 sky130_fd_sc_hd__nand2_2 _24705_ (.A(_14581_),
    .B(_14582_),
    .Y(_14583_));
 sky130_fd_sc_hd__nand2_2 _24706_ (.A(_14490_),
    .B(_14492_),
    .Y(_14584_));
 sky130_fd_sc_hd__xnor2_2 _24707_ (.A(_14583_),
    .B(_14584_),
    .Y(_14585_));
 sky130_fd_sc_hd__xnor2_2 _24708_ (.A(_14513_),
    .B(_14585_),
    .Y(_14586_));
 sky130_fd_sc_hd__nor2_2 _24709_ (.A(_14338_),
    .B(_14424_),
    .Y(_14587_));
 sky130_fd_sc_hd__a21oi_2 _24710_ (.A1(_14425_),
    .A2(_14426_),
    .B1(_14587_),
    .Y(_14588_));
 sky130_fd_sc_hd__nand2_2 _24711_ (.A(_14339_),
    .B(_14423_),
    .Y(_14589_));
 sky130_fd_sc_hd__nor2_2 _24712_ (.A(_14420_),
    .B(_14421_),
    .Y(_14590_));
 sky130_fd_sc_hd__buf_6 _24713_ (.A(_11374_),
    .X(_14592_));
 sky130_fd_sc_hd__buf_1 _24714_ (.A(_14411_),
    .X(_14593_));
 sky130_fd_sc_hd__nor2_2 _24715_ (.A(_14394_),
    .B(_14396_),
    .Y(_14594_));
 sky130_fd_sc_hd__a31o_2 _24716_ (.A1(_14592_),
    .A2(_14397_),
    .A3(_14593_),
    .B1(_14594_),
    .X(_14595_));
 sky130_fd_sc_hd__or2b_2 _24717_ (.A(_14349_),
    .B_N(_14341_),
    .X(_14596_));
 sky130_fd_sc_hd__a21bo_2 _24718_ (.A1(_14342_),
    .A2(_14348_),
    .B1_N(_14596_),
    .X(_14597_));
 sky130_fd_sc_hd__nand2_2 _24719_ (.A(iY[13]),
    .B(iY[45]),
    .Y(_14598_));
 sky130_fd_sc_hd__or2_2 _24720_ (.A(iY[13]),
    .B(iY[45]),
    .X(_14599_));
 sky130_fd_sc_hd__nand2_2 _24721_ (.A(_14598_),
    .B(_14599_),
    .Y(_14600_));
 sky130_fd_sc_hd__and3_2 _24722_ (.A(_14403_),
    .B(_14407_),
    .C(_14600_),
    .X(_14601_));
 sky130_fd_sc_hd__a21oi_2 _24723_ (.A1(_14403_),
    .A2(_14407_),
    .B1(_14600_),
    .Y(_14603_));
 sky130_fd_sc_hd__nor2_2 _24724_ (.A(_14601_),
    .B(_14603_),
    .Y(_14604_));
 sky130_fd_sc_hd__buf_1 _24725_ (.A(_14604_),
    .X(_14605_));
 sky130_fd_sc_hd__buf_1 _24726_ (.A(_14605_),
    .X(_14606_));
 sky130_fd_sc_hd__a22o_2 _24727_ (.A1(_12838_),
    .A2(_14411_),
    .B1(_14606_),
    .B2(_11374_),
    .X(_14607_));
 sky130_fd_sc_hd__buf_1 _24728_ (.A(_14604_),
    .X(_14608_));
 sky130_fd_sc_hd__nand2_2 _24729_ (.A(_12838_),
    .B(_14608_),
    .Y(_14609_));
 sky130_fd_sc_hd__or2_2 _24730_ (.A(_14412_),
    .B(_14609_),
    .X(_14610_));
 sky130_fd_sc_hd__and2_2 _24731_ (.A(_14607_),
    .B(_14610_),
    .X(_14611_));
 sky130_fd_sc_hd__buf_1 _24732_ (.A(_14386_),
    .X(_14612_));
 sky130_fd_sc_hd__or4_2 _24733_ (.A(_11827_),
    .B(_12223_),
    .C(_14612_),
    .D(_13893_),
    .X(_14614_));
 sky130_fd_sc_hd__a22o_2 _24734_ (.A1(_12225_),
    .A2(_13543_),
    .B1(_13888_),
    .B2(_14388_),
    .X(_14615_));
 sky130_fd_sc_hd__nand2_2 _24735_ (.A(_14614_),
    .B(_14615_),
    .Y(_14616_));
 sky130_fd_sc_hd__nand2_2 _24736_ (.A(_12827_),
    .B(_14392_),
    .Y(_14617_));
 sky130_fd_sc_hd__xnor2_2 _24737_ (.A(_14616_),
    .B(_14617_),
    .Y(_14618_));
 sky130_fd_sc_hd__o21a_2 _24738_ (.A1(_14390_),
    .A2(_14393_),
    .B1(_14387_),
    .X(_14619_));
 sky130_fd_sc_hd__xor2_2 _24739_ (.A(_14618_),
    .B(_14619_),
    .X(_14620_));
 sky130_fd_sc_hd__xnor2_2 _24740_ (.A(_14611_),
    .B(_14620_),
    .Y(_14621_));
 sky130_fd_sc_hd__xor2_2 _24741_ (.A(_14597_),
    .B(_14621_),
    .X(_14622_));
 sky130_fd_sc_hd__xnor2_2 _24742_ (.A(_14595_),
    .B(_14622_),
    .Y(_14623_));
 sky130_fd_sc_hd__buf_1 _24743_ (.A(_13273_),
    .X(_14625_));
 sky130_fd_sc_hd__buf_1 _24744_ (.A(_14625_),
    .X(_14626_));
 sky130_fd_sc_hd__nor2_2 _24745_ (.A(_14626_),
    .B(_14345_),
    .Y(_14627_));
 sky130_fd_sc_hd__buf_6 _24746_ (.A(_12225_),
    .X(_14628_));
 sky130_fd_sc_hd__buf_1 _24747_ (.A(_14628_),
    .X(_14629_));
 sky130_fd_sc_hd__a22o_2 _24748_ (.A1(_13953_),
    .A2(_14344_),
    .B1(_14627_),
    .B2(_14629_),
    .X(_14630_));
 sky130_fd_sc_hd__a21bo_2 _24749_ (.A1(_14354_),
    .A2(_14358_),
    .B1_N(_14353_),
    .X(_14631_));
 sky130_fd_sc_hd__nor2_2 _24750_ (.A(_12808_),
    .B(_12850_),
    .Y(_14632_));
 sky130_fd_sc_hd__nand2_2 _24751_ (.A(_14344_),
    .B(_14632_),
    .Y(_14633_));
 sky130_fd_sc_hd__inv_2 _24752_ (.A(_12772_),
    .Y(_14634_));
 sky130_fd_sc_hd__buf_1 _24753_ (.A(_14634_),
    .X(_14636_));
 sky130_fd_sc_hd__buf_1 _24754_ (.A(_12845_),
    .X(_14637_));
 sky130_fd_sc_hd__a22o_2 _24755_ (.A1(_14636_),
    .A2(_13501_),
    .B1(_14637_),
    .B2(_12816_),
    .X(_14638_));
 sky130_fd_sc_hd__nand2_2 _24756_ (.A(_14633_),
    .B(_14638_),
    .Y(_14639_));
 sky130_fd_sc_hd__buf_6 _24757_ (.A(_12457_),
    .X(_14640_));
 sky130_fd_sc_hd__buf_1 _24758_ (.A(_13273_),
    .X(_14641_));
 sky130_fd_sc_hd__or2_2 _24759_ (.A(_14640_),
    .B(_14641_),
    .X(_14642_));
 sky130_fd_sc_hd__xnor2_2 _24760_ (.A(_14639_),
    .B(_14642_),
    .Y(_14643_));
 sky130_fd_sc_hd__xor2_2 _24761_ (.A(_14631_),
    .B(_14643_),
    .X(_14644_));
 sky130_fd_sc_hd__xnor2_2 _24762_ (.A(_14630_),
    .B(_14644_),
    .Y(_14645_));
 sky130_fd_sc_hd__or4_2 _24763_ (.A(_13926_),
    .B(_12248_),
    .C(_13502_),
    .D(_13842_),
    .X(_14647_));
 sky130_fd_sc_hd__buf_1 _24764_ (.A(_13496_),
    .X(_14648_));
 sky130_fd_sc_hd__buf_1 _24765_ (.A(_11842_),
    .X(_14649_));
 sky130_fd_sc_hd__a22o_2 _24766_ (.A1(_12243_),
    .A2(_14648_),
    .B1(_13845_),
    .B2(_14649_),
    .X(_14650_));
 sky130_fd_sc_hd__nand2_2 _24767_ (.A(_14647_),
    .B(_14650_),
    .Y(_14651_));
 sky130_fd_sc_hd__buf_1 _24768_ (.A(_13244_),
    .X(_14652_));
 sky130_fd_sc_hd__nand2_2 _24769_ (.A(_12759_),
    .B(_14652_),
    .Y(_14653_));
 sky130_fd_sc_hd__xor2_2 _24770_ (.A(_14651_),
    .B(_14653_),
    .X(_14654_));
 sky130_fd_sc_hd__nand2_2 _24771_ (.A(_12451_),
    .B(_13938_),
    .Y(_14655_));
 sky130_fd_sc_hd__xnor2_2 _24772_ (.A(iX[13]),
    .B(iX[45]),
    .Y(_14656_));
 sky130_fd_sc_hd__nand2_2 _24773_ (.A(iX[12]),
    .B(iX[44]),
    .Y(_14658_));
 sky130_fd_sc_hd__o311a_2 _24774_ (.A1(_14363_),
    .A2(_14364_),
    .A3(_14366_),
    .B1(_14656_),
    .C1(_14658_),
    .X(_14659_));
 sky130_fd_sc_hd__nor2_2 _24775_ (.A(_14658_),
    .B(_14656_),
    .Y(_14660_));
 sky130_fd_sc_hd__nor2_2 _24776_ (.A(_14364_),
    .B(_14656_),
    .Y(_14661_));
 sky130_fd_sc_hd__nor3b_2 _24777_ (.A(_14363_),
    .B(_14366_),
    .C_N(_14661_),
    .Y(_14662_));
 sky130_fd_sc_hd__or4_2 _24778_ (.A(_11565_),
    .B(_14659_),
    .C(_14660_),
    .D(_14662_),
    .X(_14663_));
 sky130_fd_sc_hd__xor2_2 _24779_ (.A(_14369_),
    .B(_14663_),
    .X(_14664_));
 sky130_fd_sc_hd__xor2_2 _24780_ (.A(_14655_),
    .B(_14664_),
    .X(_14665_));
 sky130_fd_sc_hd__a22o_2 _24781_ (.A1(_14361_),
    .A2(_14369_),
    .B1(_14370_),
    .B2(_14360_),
    .X(_14666_));
 sky130_fd_sc_hd__xor2_2 _24782_ (.A(_14665_),
    .B(_14666_),
    .X(_14667_));
 sky130_fd_sc_hd__xnor2_2 _24783_ (.A(_14654_),
    .B(_14667_),
    .Y(_14669_));
 sky130_fd_sc_hd__nor2_2 _24784_ (.A(_14372_),
    .B(_14374_),
    .Y(_14670_));
 sky130_fd_sc_hd__a21o_2 _24785_ (.A1(_14359_),
    .A2(_14375_),
    .B1(_14670_),
    .X(_14671_));
 sky130_fd_sc_hd__xnor2_2 _24786_ (.A(_14669_),
    .B(_14671_),
    .Y(_14672_));
 sky130_fd_sc_hd__xnor2_2 _24787_ (.A(_14645_),
    .B(_14672_),
    .Y(_14673_));
 sky130_fd_sc_hd__nor2_2 _24788_ (.A(_14376_),
    .B(_14377_),
    .Y(_14674_));
 sky130_fd_sc_hd__a21o_2 _24789_ (.A1(_14350_),
    .A2(_14378_),
    .B1(_14674_),
    .X(_14675_));
 sky130_fd_sc_hd__xnor2_2 _24790_ (.A(_14673_),
    .B(_14675_),
    .Y(_14676_));
 sky130_fd_sc_hd__xnor2_2 _24791_ (.A(_14623_),
    .B(_14676_),
    .Y(_14677_));
 sky130_fd_sc_hd__nor2_2 _24792_ (.A(_14379_),
    .B(_14380_),
    .Y(_14678_));
 sky130_fd_sc_hd__a21oi_2 _24793_ (.A1(_14381_),
    .A2(_14415_),
    .B1(_14678_),
    .Y(_14680_));
 sky130_fd_sc_hd__xnor2_2 _24794_ (.A(_14677_),
    .B(_14680_),
    .Y(_14681_));
 sky130_fd_sc_hd__nand2_2 _24795_ (.A(_14385_),
    .B(_14413_),
    .Y(_14682_));
 sky130_fd_sc_hd__o21ai_2 _24796_ (.A1(_14382_),
    .A2(_14414_),
    .B1(_14682_),
    .Y(_14683_));
 sky130_fd_sc_hd__xor2_2 _24797_ (.A(_14681_),
    .B(_14683_),
    .X(_14684_));
 sky130_fd_sc_hd__and2b_2 _24798_ (.A_N(_14418_),
    .B(_14416_),
    .X(_14685_));
 sky130_fd_sc_hd__a21o_2 _24799_ (.A1(_13976_),
    .A2(_14419_),
    .B1(_14685_),
    .X(_14686_));
 sky130_fd_sc_hd__xor2_2 _24800_ (.A(_14684_),
    .B(_14686_),
    .X(_14687_));
 sky130_fd_sc_hd__xor2_2 _24801_ (.A(_14590_),
    .B(_14687_),
    .X(_14688_));
 sky130_fd_sc_hd__or3_4 _24802_ (.A(_14336_),
    .B(_14422_),
    .C(_14688_),
    .X(_14689_));
 sky130_fd_sc_hd__o21ai_2 _24803_ (.A1(_14336_),
    .A2(_14422_),
    .B1(_14688_),
    .Y(_14691_));
 sky130_fd_sc_hd__a21bo_2 _24804_ (.A1(_14689_),
    .A2(_14691_),
    .B1_N(_14589_),
    .X(_14692_));
 sky130_fd_sc_hd__o21a_2 _24805_ (.A1(_14589_),
    .A2(_14688_),
    .B1(_14692_),
    .X(_14693_));
 sky130_fd_sc_hd__xnor2_2 _24806_ (.A(_14588_),
    .B(_14693_),
    .Y(_14694_));
 sky130_fd_sc_hd__xor2_2 _24807_ (.A(_14586_),
    .B(_14694_),
    .X(_14695_));
 sky130_fd_sc_hd__xor2_2 _24808_ (.A(oO[13]),
    .B(_14695_),
    .X(_14696_));
 sky130_fd_sc_hd__and2b_2 _24809_ (.A_N(oO[12]),
    .B(_14500_),
    .X(_14697_));
 sky130_fd_sc_hd__a21oi_2 _24810_ (.A1(_14427_),
    .A2(_14499_),
    .B1(_14697_),
    .Y(_14698_));
 sky130_fd_sc_hd__xnor2_2 _24811_ (.A(_14696_),
    .B(_14698_),
    .Y(_14699_));
 sky130_fd_sc_hd__nor2_2 _24812_ (.A(_14501_),
    .B(_14502_),
    .Y(_14700_));
 sky130_fd_sc_hd__a21oi_2 _24813_ (.A1(_14503_),
    .A2(_14506_),
    .B1(_14700_),
    .Y(_14702_));
 sky130_fd_sc_hd__xor2_2 _24814_ (.A(_14699_),
    .B(_14702_),
    .X(_14703_));
 sky130_fd_sc_hd__and2b_2 _24815_ (.A_N(_14315_),
    .B(_14316_),
    .X(_14704_));
 sky130_fd_sc_hd__nand2_2 _24816_ (.A(iY[14]),
    .B(iX[31]),
    .Y(_14705_));
 sky130_fd_sc_hd__a21o_2 _24817_ (.A1(_14118_),
    .A2(_14233_),
    .B1(_14244_),
    .X(_14706_));
 sky130_fd_sc_hd__nand2_2 _24818_ (.A(_14234_),
    .B(_14243_),
    .Y(_14707_));
 sky130_fd_sc_hd__and2_2 _24819_ (.A(iY[16]),
    .B(iX[30]),
    .X(_14708_));
 sky130_fd_sc_hd__and3_2 _24820_ (.A(iY[15]),
    .B(iX[29]),
    .C(_14708_),
    .X(_14709_));
 sky130_fd_sc_hd__a22oi_2 _24821_ (.A1(iY[16]),
    .A2(iX[29]),
    .B1(iX[30]),
    .B2(iY[15]),
    .Y(_14710_));
 sky130_fd_sc_hd__nor2_2 _24822_ (.A(_14709_),
    .B(_14710_),
    .Y(_14711_));
 sky130_fd_sc_hd__nand2_2 _24823_ (.A(iY[17]),
    .B(iX[28]),
    .Y(_14713_));
 sky130_fd_sc_hd__xnor2_2 _24824_ (.A(_14711_),
    .B(_14713_),
    .Y(_14714_));
 sky130_fd_sc_hd__and2_2 _24825_ (.A(_14214_),
    .B(_14714_),
    .X(_14715_));
 sky130_fd_sc_hd__nor2_2 _24826_ (.A(_14214_),
    .B(_14714_),
    .Y(_14716_));
 sky130_fd_sc_hd__or2_2 _24827_ (.A(_14715_),
    .B(_14716_),
    .X(_14717_));
 sky130_fd_sc_hd__a31o_2 _24828_ (.A1(iY[17]),
    .A2(iX[27]),
    .A3(_14237_),
    .B1(_14235_),
    .X(_14718_));
 sky130_fd_sc_hd__and2b_2 _24829_ (.A_N(_14717_),
    .B(_14718_),
    .X(_14719_));
 sky130_fd_sc_hd__and2b_2 _24830_ (.A_N(_14718_),
    .B(_14717_),
    .X(_14720_));
 sky130_fd_sc_hd__or2_2 _24831_ (.A(_14719_),
    .B(_14720_),
    .X(_14721_));
 sky130_fd_sc_hd__a21oi_2 _24832_ (.A1(_14240_),
    .A2(_14707_),
    .B1(_14721_),
    .Y(_14722_));
 sky130_fd_sc_hd__and3_2 _24833_ (.A(_14240_),
    .B(_14707_),
    .C(_14721_),
    .X(_14724_));
 sky130_fd_sc_hd__and4_2 _24834_ (.A(iY[21]),
    .B(iY[22]),
    .C(iX[23]),
    .D(iX[24]),
    .X(_14725_));
 sky130_fd_sc_hd__a22oi_2 _24835_ (.A1(iY[22]),
    .A2(iX[23]),
    .B1(iX[24]),
    .B2(iY[21]),
    .Y(_14726_));
 sky130_fd_sc_hd__nor2_2 _24836_ (.A(_14725_),
    .B(_14726_),
    .Y(_14727_));
 sky130_fd_sc_hd__nand2_2 _24837_ (.A(iX[22]),
    .B(iY[23]),
    .Y(_14728_));
 sky130_fd_sc_hd__xnor2_2 _24838_ (.A(_14727_),
    .B(_14728_),
    .Y(_14729_));
 sky130_fd_sc_hd__and4_2 _24839_ (.A(iY[18]),
    .B(iY[19]),
    .C(iX[26]),
    .D(iX[27]),
    .X(_14730_));
 sky130_fd_sc_hd__a22oi_2 _24840_ (.A1(iY[19]),
    .A2(iX[26]),
    .B1(iX[27]),
    .B2(iY[18]),
    .Y(_14731_));
 sky130_fd_sc_hd__nor2_2 _24841_ (.A(_14730_),
    .B(_14731_),
    .Y(_14732_));
 sky130_fd_sc_hd__nand2_2 _24842_ (.A(iY[20]),
    .B(iX[25]),
    .Y(_14733_));
 sky130_fd_sc_hd__xnor2_2 _24843_ (.A(_14732_),
    .B(_14733_),
    .Y(_14735_));
 sky130_fd_sc_hd__o21ba_2 _24844_ (.A1(_14223_),
    .A2(_14225_),
    .B1_N(_14222_),
    .X(_14736_));
 sky130_fd_sc_hd__xnor2_2 _24845_ (.A(_14735_),
    .B(_14736_),
    .Y(_14737_));
 sky130_fd_sc_hd__and2_2 _24846_ (.A(_14729_),
    .B(_14737_),
    .X(_14738_));
 sky130_fd_sc_hd__nor2_2 _24847_ (.A(_14729_),
    .B(_14737_),
    .Y(_14739_));
 sky130_fd_sc_hd__or2_2 _24848_ (.A(_14738_),
    .B(_14739_),
    .X(_14740_));
 sky130_fd_sc_hd__nor3_2 _24849_ (.A(_14722_),
    .B(_14724_),
    .C(_14740_),
    .Y(_14741_));
 sky130_fd_sc_hd__o21a_2 _24850_ (.A1(_14722_),
    .A2(_14724_),
    .B1(_14740_),
    .X(_14742_));
 sky130_fd_sc_hd__a211oi_2 _24851_ (.A1(_14706_),
    .A2(_14247_),
    .B1(_14741_),
    .C1(_14742_),
    .Y(_14743_));
 sky130_fd_sc_hd__o211a_2 _24852_ (.A1(_14741_),
    .A2(_14742_),
    .B1(_14706_),
    .C1(_14247_),
    .X(_14744_));
 sky130_fd_sc_hd__nor2_2 _24853_ (.A(_14743_),
    .B(_14744_),
    .Y(_14746_));
 sky130_fd_sc_hd__xnor2_2 _24854_ (.A(_14705_),
    .B(_14746_),
    .Y(_14747_));
 sky130_fd_sc_hd__xnor2_2 _24855_ (.A(_14254_),
    .B(_14747_),
    .Y(_14748_));
 sky130_fd_sc_hd__inv_2 _24856_ (.A(_14300_),
    .Y(_14749_));
 sky130_fd_sc_hd__or2b_2 _24857_ (.A(_14268_),
    .B_N(_14267_),
    .X(_14750_));
 sky130_fd_sc_hd__and4_2 _24858_ (.A(iX[17]),
    .B(iX[18]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_14751_));
 sky130_fd_sc_hd__a22oi_2 _24859_ (.A1(iX[18]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[17]),
    .Y(_14752_));
 sky130_fd_sc_hd__nor2_2 _24860_ (.A(_14751_),
    .B(_14752_),
    .Y(_14753_));
 sky130_fd_sc_hd__nand2_2 _24861_ (.A(iX[16]),
    .B(iY[29]),
    .Y(_14754_));
 sky130_fd_sc_hd__xnor2_2 _24862_ (.A(_14753_),
    .B(_14754_),
    .Y(_14755_));
 sky130_fd_sc_hd__o21ba_2 _24863_ (.A1(_14264_),
    .A2(_14266_),
    .B1_N(_14262_),
    .X(_14757_));
 sky130_fd_sc_hd__xnor2_2 _24864_ (.A(_14755_),
    .B(_14757_),
    .Y(_14758_));
 sky130_fd_sc_hd__nand3_2 _24865_ (.A(iX[15]),
    .B(iY[30]),
    .C(_14758_),
    .Y(_14759_));
 sky130_fd_sc_hd__a21o_2 _24866_ (.A1(iX[15]),
    .A2(iY[30]),
    .B1(_14758_),
    .X(_14760_));
 sky130_fd_sc_hd__nand2_2 _24867_ (.A(_14759_),
    .B(_14760_),
    .Y(_14761_));
 sky130_fd_sc_hd__a21oi_2 _24868_ (.A1(_14750_),
    .A2(_14270_),
    .B1(_14761_),
    .Y(_14762_));
 sky130_fd_sc_hd__and3_2 _24869_ (.A(_14750_),
    .B(_14270_),
    .C(_14761_),
    .X(_14763_));
 sky130_fd_sc_hd__nor2_2 _24870_ (.A(_14762_),
    .B(_14763_),
    .Y(_14764_));
 sky130_fd_sc_hd__a21oi_2 _24871_ (.A1(iX[14]),
    .A2(iY[31]),
    .B1(_14764_),
    .Y(_14765_));
 sky130_fd_sc_hd__and3_2 _24872_ (.A(iX[14]),
    .B(iY[31]),
    .C(_14764_),
    .X(_14766_));
 sky130_fd_sc_hd__nor2_2 _24873_ (.A(_14765_),
    .B(_14766_),
    .Y(_14768_));
 sky130_fd_sc_hd__or2b_2 _24874_ (.A(_14286_),
    .B_N(_14291_),
    .X(_14769_));
 sky130_fd_sc_hd__or2b_2 _24875_ (.A(_14284_),
    .B_N(_14292_),
    .X(_14770_));
 sky130_fd_sc_hd__and2b_2 _24876_ (.A_N(_14227_),
    .B(_14226_),
    .X(_14771_));
 sky130_fd_sc_hd__o21ba_2 _24877_ (.A1(_14288_),
    .A2(_14290_),
    .B1_N(_14287_),
    .X(_14772_));
 sky130_fd_sc_hd__o21ba_2 _24878_ (.A1(_14217_),
    .A2(_14220_),
    .B1_N(_14216_),
    .X(_14773_));
 sky130_fd_sc_hd__and4_2 _24879_ (.A(iX[20]),
    .B(iX[21]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_14774_));
 sky130_fd_sc_hd__a22oi_2 _24880_ (.A1(iX[21]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[20]),
    .Y(_14775_));
 sky130_fd_sc_hd__nor2_2 _24881_ (.A(_14774_),
    .B(_14775_),
    .Y(_14776_));
 sky130_fd_sc_hd__nand2_2 _24882_ (.A(iX[19]),
    .B(iY[26]),
    .Y(_14777_));
 sky130_fd_sc_hd__xnor2_2 _24883_ (.A(_14776_),
    .B(_14777_),
    .Y(_14779_));
 sky130_fd_sc_hd__xnor2_2 _24884_ (.A(_14773_),
    .B(_14779_),
    .Y(_14780_));
 sky130_fd_sc_hd__xnor2_2 _24885_ (.A(_14772_),
    .B(_14780_),
    .Y(_14781_));
 sky130_fd_sc_hd__o21a_2 _24886_ (.A1(_14771_),
    .A2(_14229_),
    .B1(_14781_),
    .X(_14782_));
 sky130_fd_sc_hd__nor3_2 _24887_ (.A(_14771_),
    .B(_14229_),
    .C(_14781_),
    .Y(_14783_));
 sky130_fd_sc_hd__a211oi_2 _24888_ (.A1(_14769_),
    .A2(_14770_),
    .B1(_14782_),
    .C1(_14783_),
    .Y(_14784_));
 sky130_fd_sc_hd__o211a_2 _24889_ (.A1(_14782_),
    .A2(_14783_),
    .B1(_14769_),
    .C1(_14770_),
    .X(_14785_));
 sky130_fd_sc_hd__nor2_2 _24890_ (.A(_14294_),
    .B(_14297_),
    .Y(_14786_));
 sky130_fd_sc_hd__or3_2 _24891_ (.A(_14784_),
    .B(_14785_),
    .C(_14786_),
    .X(_14787_));
 sky130_fd_sc_hd__o21ai_2 _24892_ (.A1(_14784_),
    .A2(_14785_),
    .B1(_14786_),
    .Y(_14788_));
 sky130_fd_sc_hd__nand3_2 _24893_ (.A(_14768_),
    .B(_14787_),
    .C(_14788_),
    .Y(_14790_));
 sky130_fd_sc_hd__a21o_2 _24894_ (.A1(_14787_),
    .A2(_14788_),
    .B1(_14768_),
    .X(_14791_));
 sky130_fd_sc_hd__and2_2 _24895_ (.A(_14790_),
    .B(_14791_),
    .X(_14792_));
 sky130_fd_sc_hd__o21ai_2 _24896_ (.A1(_14249_),
    .A2(_14251_),
    .B1(_14792_),
    .Y(_14793_));
 sky130_fd_sc_hd__or3_2 _24897_ (.A(_14249_),
    .B(_14251_),
    .C(_14792_),
    .X(_14794_));
 sky130_fd_sc_hd__o211ai_2 _24898_ (.A1(_14749_),
    .A2(_14302_),
    .B1(_14793_),
    .C1(_14794_),
    .Y(_14795_));
 sky130_fd_sc_hd__a211o_2 _24899_ (.A1(_14793_),
    .A2(_14794_),
    .B1(_14749_),
    .C1(_14302_),
    .X(_14796_));
 sky130_fd_sc_hd__and3_2 _24900_ (.A(_14748_),
    .B(_14795_),
    .C(_14796_),
    .X(_14797_));
 sky130_fd_sc_hd__a21oi_2 _24901_ (.A1(_14795_),
    .A2(_14796_),
    .B1(_14748_),
    .Y(_14798_));
 sky130_fd_sc_hd__a211oi_2 _24902_ (.A1(_14256_),
    .A2(_14310_),
    .B1(_14797_),
    .C1(_14798_),
    .Y(_14799_));
 sky130_fd_sc_hd__o211a_2 _24903_ (.A1(_14797_),
    .A2(_14798_),
    .B1(_14256_),
    .C1(_14310_),
    .X(_14801_));
 sky130_fd_sc_hd__a211oi_2 _24904_ (.A1(_14304_),
    .A2(_14308_),
    .B1(_14799_),
    .C1(_14801_),
    .Y(_14802_));
 sky130_fd_sc_hd__o211a_2 _24905_ (.A1(_14799_),
    .A2(_14801_),
    .B1(_14304_),
    .C1(_14308_),
    .X(_14803_));
 sky130_fd_sc_hd__nor2_2 _24906_ (.A(_14802_),
    .B(_14803_),
    .Y(_14804_));
 sky130_fd_sc_hd__o21a_2 _24907_ (.A1(_14313_),
    .A2(_14704_),
    .B1(_14804_),
    .X(_14805_));
 sky130_fd_sc_hd__nor3_2 _24908_ (.A(_14313_),
    .B(_14704_),
    .C(_14804_),
    .Y(_14806_));
 sky130_fd_sc_hd__a211oi_2 _24909_ (.A1(_14273_),
    .A2(_14279_),
    .B1(_14805_),
    .C1(_14806_),
    .Y(_14807_));
 sky130_fd_sc_hd__o211a_2 _24910_ (.A1(_14805_),
    .A2(_14806_),
    .B1(_14273_),
    .C1(_14279_),
    .X(_14808_));
 sky130_fd_sc_hd__a211o_2 _24911_ (.A1(_14319_),
    .A2(_14322_),
    .B1(_14807_),
    .C1(_14808_),
    .X(_14809_));
 sky130_fd_sc_hd__inv_2 _24912_ (.A(_14809_),
    .Y(_14810_));
 sky130_fd_sc_hd__o211a_2 _24913_ (.A1(_14807_),
    .A2(_14808_),
    .B1(_14319_),
    .C1(_14322_),
    .X(_14812_));
 sky130_fd_sc_hd__nor2_2 _24914_ (.A(_14810_),
    .B(_14812_),
    .Y(_14813_));
 sky130_fd_sc_hd__nor2_2 _24915_ (.A(_14326_),
    .B(_14330_),
    .Y(_14814_));
 sky130_fd_sc_hd__xnor2_2 _24916_ (.A(_14813_),
    .B(_14814_),
    .Y(_14815_));
 sky130_fd_sc_hd__nand2_2 _24917_ (.A(_14703_),
    .B(_14815_),
    .Y(_14816_));
 sky130_fd_sc_hd__nor2_2 _24918_ (.A(_14703_),
    .B(_14815_),
    .Y(_14817_));
 sky130_fd_sc_hd__inv_2 _24919_ (.A(_14817_),
    .Y(_14818_));
 sky130_fd_sc_hd__nand2_2 _24920_ (.A(_14816_),
    .B(_14818_),
    .Y(_14819_));
 sky130_fd_sc_hd__and2b_2 _24921_ (.A_N(_14335_),
    .B(_14507_),
    .X(_14820_));
 sky130_fd_sc_hd__or2_2 _24922_ (.A(_14820_),
    .B(_14510_),
    .X(_14821_));
 sky130_fd_sc_hd__xnor2_2 _24923_ (.A(_14819_),
    .B(_14821_),
    .Y(oO[45]));
 sky130_fd_sc_hd__and2b_2 _24924_ (.A_N(_14254_),
    .B(_14747_),
    .X(_14823_));
 sky130_fd_sc_hd__or3_2 _24925_ (.A(_14705_),
    .B(_14743_),
    .C(_14744_),
    .X(_14824_));
 sky130_fd_sc_hd__and3_2 _24926_ (.A(iY[15]),
    .B(iX[31]),
    .C(_14708_),
    .X(_14825_));
 sky130_fd_sc_hd__a21o_2 _24927_ (.A1(iY[15]),
    .A2(iX[31]),
    .B1(_14708_),
    .X(_14826_));
 sky130_fd_sc_hd__and2b_2 _24928_ (.A_N(_14825_),
    .B(_14826_),
    .X(_14827_));
 sky130_fd_sc_hd__nand2_2 _24929_ (.A(iY[17]),
    .B(iX[29]),
    .Y(_14828_));
 sky130_fd_sc_hd__xnor2_2 _24930_ (.A(_14827_),
    .B(_14828_),
    .Y(_14829_));
 sky130_fd_sc_hd__o21ba_2 _24931_ (.A1(_14710_),
    .A2(_14713_),
    .B1_N(_14709_),
    .X(_14830_));
 sky130_fd_sc_hd__xnor2_2 _24932_ (.A(_14829_),
    .B(_14830_),
    .Y(_14831_));
 sky130_fd_sc_hd__o21a_2 _24933_ (.A1(_14715_),
    .A2(_14719_),
    .B1(_14831_),
    .X(_14833_));
 sky130_fd_sc_hd__nor3_2 _24934_ (.A(_14715_),
    .B(_14719_),
    .C(_14831_),
    .Y(_14834_));
 sky130_fd_sc_hd__nor2_2 _24935_ (.A(_14833_),
    .B(_14834_),
    .Y(_14835_));
 sky130_fd_sc_hd__and4_2 _24936_ (.A(iY[21]),
    .B(iY[22]),
    .C(iX[24]),
    .D(iX[25]),
    .X(_14836_));
 sky130_fd_sc_hd__a22oi_2 _24937_ (.A1(iY[22]),
    .A2(iX[24]),
    .B1(iX[25]),
    .B2(iY[21]),
    .Y(_14837_));
 sky130_fd_sc_hd__nor2_2 _24938_ (.A(_14836_),
    .B(_14837_),
    .Y(_14838_));
 sky130_fd_sc_hd__nand2_2 _24939_ (.A(iX[23]),
    .B(iY[23]),
    .Y(_14839_));
 sky130_fd_sc_hd__xnor2_2 _24940_ (.A(_14838_),
    .B(_14839_),
    .Y(_14840_));
 sky130_fd_sc_hd__and4_2 _24941_ (.A(iY[18]),
    .B(iY[19]),
    .C(iX[27]),
    .D(iX[28]),
    .X(_14841_));
 sky130_fd_sc_hd__a22oi_2 _24942_ (.A1(iY[19]),
    .A2(iX[27]),
    .B1(iX[28]),
    .B2(iY[18]),
    .Y(_14842_));
 sky130_fd_sc_hd__nor2_2 _24943_ (.A(_14841_),
    .B(_14842_),
    .Y(_14844_));
 sky130_fd_sc_hd__nand2_2 _24944_ (.A(iY[20]),
    .B(iX[26]),
    .Y(_14845_));
 sky130_fd_sc_hd__xnor2_2 _24945_ (.A(_14844_),
    .B(_14845_),
    .Y(_14846_));
 sky130_fd_sc_hd__o21ba_2 _24946_ (.A1(_14731_),
    .A2(_14733_),
    .B1_N(_14730_),
    .X(_14847_));
 sky130_fd_sc_hd__xnor2_2 _24947_ (.A(_14846_),
    .B(_14847_),
    .Y(_14848_));
 sky130_fd_sc_hd__and2_2 _24948_ (.A(_14840_),
    .B(_14848_),
    .X(_14849_));
 sky130_fd_sc_hd__nor2_2 _24949_ (.A(_14840_),
    .B(_14848_),
    .Y(_14850_));
 sky130_fd_sc_hd__or2_2 _24950_ (.A(_14849_),
    .B(_14850_),
    .X(_14851_));
 sky130_fd_sc_hd__inv_2 _24951_ (.A(_14851_),
    .Y(_14852_));
 sky130_fd_sc_hd__xnor2_2 _24952_ (.A(_14835_),
    .B(_14852_),
    .Y(_14853_));
 sky130_fd_sc_hd__o21ba_2 _24953_ (.A1(_14722_),
    .A2(_14741_),
    .B1_N(_14853_),
    .X(_14855_));
 sky130_fd_sc_hd__or3b_2 _24954_ (.A(_14722_),
    .B(_14741_),
    .C_N(_14853_),
    .X(_14856_));
 sky130_fd_sc_hd__or2b_2 _24955_ (.A(_14855_),
    .B_N(_14856_),
    .X(_14857_));
 sky130_fd_sc_hd__xnor2_2 _24956_ (.A(_14824_),
    .B(_14857_),
    .Y(_14858_));
 sky130_fd_sc_hd__or2b_2 _24957_ (.A(_14757_),
    .B_N(_14755_),
    .X(_14859_));
 sky130_fd_sc_hd__and4_2 _24958_ (.A(iX[18]),
    .B(iX[19]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_14860_));
 sky130_fd_sc_hd__a22oi_2 _24959_ (.A1(iX[19]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[18]),
    .Y(_14861_));
 sky130_fd_sc_hd__nor2_2 _24960_ (.A(_14860_),
    .B(_14861_),
    .Y(_14862_));
 sky130_fd_sc_hd__nand2_2 _24961_ (.A(iX[17]),
    .B(iY[29]),
    .Y(_14863_));
 sky130_fd_sc_hd__xnor2_2 _24962_ (.A(_14862_),
    .B(_14863_),
    .Y(_14864_));
 sky130_fd_sc_hd__o21ba_2 _24963_ (.A1(_14752_),
    .A2(_14754_),
    .B1_N(_14751_),
    .X(_14866_));
 sky130_fd_sc_hd__xnor2_2 _24964_ (.A(_14864_),
    .B(_14866_),
    .Y(_14867_));
 sky130_fd_sc_hd__and2_2 _24965_ (.A(iX[16]),
    .B(iY[30]),
    .X(_14868_));
 sky130_fd_sc_hd__or2_2 _24966_ (.A(_14867_),
    .B(_14868_),
    .X(_14869_));
 sky130_fd_sc_hd__nand2_2 _24967_ (.A(_14867_),
    .B(_14868_),
    .Y(_14870_));
 sky130_fd_sc_hd__nand2_2 _24968_ (.A(_14869_),
    .B(_14870_),
    .Y(_14871_));
 sky130_fd_sc_hd__a21oi_2 _24969_ (.A1(_14859_),
    .A2(_14759_),
    .B1(_14871_),
    .Y(_14872_));
 sky130_fd_sc_hd__and3_2 _24970_ (.A(_14859_),
    .B(_14759_),
    .C(_14871_),
    .X(_14873_));
 sky130_fd_sc_hd__nor2_2 _24971_ (.A(_14872_),
    .B(_14873_),
    .Y(_14874_));
 sky130_fd_sc_hd__nand2_2 _24972_ (.A(iX[15]),
    .B(iY[31]),
    .Y(_14875_));
 sky130_fd_sc_hd__xnor2_2 _24973_ (.A(_14874_),
    .B(_14875_),
    .Y(_14877_));
 sky130_fd_sc_hd__or2b_2 _24974_ (.A(_14773_),
    .B_N(_14779_),
    .X(_14878_));
 sky130_fd_sc_hd__or2b_2 _24975_ (.A(_14772_),
    .B_N(_14780_),
    .X(_14879_));
 sky130_fd_sc_hd__and2b_2 _24976_ (.A_N(_14736_),
    .B(_14735_),
    .X(_14880_));
 sky130_fd_sc_hd__o21ba_2 _24977_ (.A1(_14775_),
    .A2(_14777_),
    .B1_N(_14774_),
    .X(_14881_));
 sky130_fd_sc_hd__o21ba_2 _24978_ (.A1(_14726_),
    .A2(_14728_),
    .B1_N(_14725_),
    .X(_14882_));
 sky130_fd_sc_hd__and4_2 _24979_ (.A(iX[21]),
    .B(iX[22]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_14883_));
 sky130_fd_sc_hd__a22oi_2 _24980_ (.A1(iX[22]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[21]),
    .Y(_14884_));
 sky130_fd_sc_hd__nor2_2 _24981_ (.A(_14883_),
    .B(_14884_),
    .Y(_14885_));
 sky130_fd_sc_hd__nand2_2 _24982_ (.A(iX[20]),
    .B(iY[26]),
    .Y(_14886_));
 sky130_fd_sc_hd__xnor2_2 _24983_ (.A(_14885_),
    .B(_14886_),
    .Y(_14888_));
 sky130_fd_sc_hd__xnor2_2 _24984_ (.A(_14882_),
    .B(_14888_),
    .Y(_14889_));
 sky130_fd_sc_hd__xnor2_2 _24985_ (.A(_14881_),
    .B(_14889_),
    .Y(_14890_));
 sky130_fd_sc_hd__o21a_2 _24986_ (.A1(_14880_),
    .A2(_14738_),
    .B1(_14890_),
    .X(_14891_));
 sky130_fd_sc_hd__nor3_2 _24987_ (.A(_14880_),
    .B(_14738_),
    .C(_14890_),
    .Y(_14892_));
 sky130_fd_sc_hd__a211oi_2 _24988_ (.A1(_14878_),
    .A2(_14879_),
    .B1(_14891_),
    .C1(_14892_),
    .Y(_14893_));
 sky130_fd_sc_hd__o211a_2 _24989_ (.A1(_14891_),
    .A2(_14892_),
    .B1(_14878_),
    .C1(_14879_),
    .X(_14894_));
 sky130_fd_sc_hd__nor2_2 _24990_ (.A(_14782_),
    .B(_14784_),
    .Y(_14895_));
 sky130_fd_sc_hd__or3_2 _24991_ (.A(_14893_),
    .B(_14894_),
    .C(_14895_),
    .X(_14896_));
 sky130_fd_sc_hd__o21ai_2 _24992_ (.A1(_14893_),
    .A2(_14894_),
    .B1(_14895_),
    .Y(_14897_));
 sky130_fd_sc_hd__nand3_2 _24993_ (.A(_14877_),
    .B(_14896_),
    .C(_14897_),
    .Y(_14899_));
 sky130_fd_sc_hd__a21o_2 _24994_ (.A1(_14896_),
    .A2(_14897_),
    .B1(_14877_),
    .X(_14900_));
 sky130_fd_sc_hd__and3_2 _24995_ (.A(_14743_),
    .B(_14899_),
    .C(_14900_),
    .X(_14901_));
 sky130_fd_sc_hd__a21oi_2 _24996_ (.A1(_14899_),
    .A2(_14900_),
    .B1(_14743_),
    .Y(_14902_));
 sky130_fd_sc_hd__a211oi_2 _24997_ (.A1(_14787_),
    .A2(_14790_),
    .B1(_14901_),
    .C1(_14902_),
    .Y(_14903_));
 sky130_fd_sc_hd__o211a_2 _24998_ (.A1(_14901_),
    .A2(_14902_),
    .B1(_14787_),
    .C1(_14790_),
    .X(_14904_));
 sky130_fd_sc_hd__or3_2 _24999_ (.A(_14858_),
    .B(_14903_),
    .C(_14904_),
    .X(_14905_));
 sky130_fd_sc_hd__o21ai_2 _25000_ (.A1(_14903_),
    .A2(_14904_),
    .B1(_14858_),
    .Y(_14906_));
 sky130_fd_sc_hd__o211a_2 _25001_ (.A1(_14823_),
    .A2(_14797_),
    .B1(_14905_),
    .C1(_14906_),
    .X(_14907_));
 sky130_fd_sc_hd__a211oi_2 _25002_ (.A1(_14905_),
    .A2(_14906_),
    .B1(_14823_),
    .C1(_14797_),
    .Y(_14908_));
 sky130_fd_sc_hd__or2_2 _25003_ (.A(_14907_),
    .B(_14908_),
    .X(_14910_));
 sky130_fd_sc_hd__nand2_2 _25004_ (.A(_14793_),
    .B(_14795_),
    .Y(_14911_));
 sky130_fd_sc_hd__xnor2_2 _25005_ (.A(_14910_),
    .B(_14911_),
    .Y(_14912_));
 sky130_fd_sc_hd__nor2_2 _25006_ (.A(_14799_),
    .B(_14802_),
    .Y(_14913_));
 sky130_fd_sc_hd__xnor2_2 _25007_ (.A(_14912_),
    .B(_14913_),
    .Y(_14914_));
 sky130_fd_sc_hd__o21a_2 _25008_ (.A1(_14762_),
    .A2(_14766_),
    .B1(_14914_),
    .X(_14915_));
 sky130_fd_sc_hd__nor3_2 _25009_ (.A(_14762_),
    .B(_14766_),
    .C(_14914_),
    .Y(_14916_));
 sky130_fd_sc_hd__or2_2 _25010_ (.A(_14915_),
    .B(_14916_),
    .X(_14917_));
 sky130_fd_sc_hd__nor2_2 _25011_ (.A(_14805_),
    .B(_14807_),
    .Y(_14918_));
 sky130_fd_sc_hd__nor2_2 _25012_ (.A(_14917_),
    .B(_14918_),
    .Y(_14919_));
 sky130_fd_sc_hd__and2_2 _25013_ (.A(_14917_),
    .B(_14918_),
    .X(_14921_));
 sky130_fd_sc_hd__nor2_2 _25014_ (.A(_14919_),
    .B(_14921_),
    .Y(_14922_));
 sky130_fd_sc_hd__o21bai_2 _25015_ (.A1(_14326_),
    .A2(_14810_),
    .B1_N(_14812_),
    .Y(_14923_));
 sky130_fd_sc_hd__a21bo_2 _25016_ (.A1(_14330_),
    .A2(_14813_),
    .B1_N(_14923_),
    .X(_14924_));
 sky130_fd_sc_hd__xnor2_2 _25017_ (.A(_14922_),
    .B(_14924_),
    .Y(_14925_));
 sky130_fd_sc_hd__or3_2 _25018_ (.A(_14420_),
    .B(_14421_),
    .C(_14687_),
    .X(_14926_));
 sky130_fd_sc_hd__and2b_2 _25019_ (.A_N(_14684_),
    .B(_14686_),
    .X(_14927_));
 sky130_fd_sc_hd__and2b_2 _25020_ (.A_N(_14621_),
    .B(_14597_),
    .X(_14928_));
 sky130_fd_sc_hd__and2b_2 _25021_ (.A_N(_14622_),
    .B(_14595_),
    .X(_14929_));
 sky130_fd_sc_hd__nor2_2 _25022_ (.A(_14928_),
    .B(_14929_),
    .Y(_14930_));
 sky130_fd_sc_hd__nor2_2 _25023_ (.A(_14610_),
    .B(_14930_),
    .Y(_14932_));
 sky130_fd_sc_hd__and2_2 _25024_ (.A(_14610_),
    .B(_14930_),
    .X(_14933_));
 sky130_fd_sc_hd__nor2_2 _25025_ (.A(_14932_),
    .B(_14933_),
    .Y(_14934_));
 sky130_fd_sc_hd__a2bb2o_2 _25026_ (.A1_N(_14618_),
    .A2_N(_14619_),
    .B1(_14620_),
    .B2(_14611_),
    .X(_14935_));
 sky130_fd_sc_hd__and2b_2 _25027_ (.A_N(_14643_),
    .B(_14631_),
    .X(_14936_));
 sky130_fd_sc_hd__and2b_2 _25028_ (.A_N(_14644_),
    .B(_14630_),
    .X(_14937_));
 sky130_fd_sc_hd__nand2_2 _25029_ (.A(_12827_),
    .B(_14409_),
    .Y(_14938_));
 sky130_fd_sc_hd__xor2_2 _25030_ (.A(_14609_),
    .B(_14938_),
    .X(_14939_));
 sky130_fd_sc_hd__and2_2 _25031_ (.A(iY[14]),
    .B(iY[46]),
    .X(_14940_));
 sky130_fd_sc_hd__nor2_2 _25032_ (.A(iY[14]),
    .B(iY[46]),
    .Y(_14941_));
 sky130_fd_sc_hd__nor2_2 _25033_ (.A(_14940_),
    .B(_14941_),
    .Y(_14943_));
 sky130_fd_sc_hd__nor2_2 _25034_ (.A(_14405_),
    .B(_14600_),
    .Y(_14944_));
 sky130_fd_sc_hd__nand2_2 _25035_ (.A(_14403_),
    .B(_14598_),
    .Y(_14945_));
 sky130_fd_sc_hd__a22o_2 _25036_ (.A1(_14599_),
    .A2(_14945_),
    .B1(_14944_),
    .B2(_14400_),
    .X(_14946_));
 sky130_fd_sc_hd__a21o_4 _25037_ (.A1(_14402_),
    .A2(_14944_),
    .B1(_14946_),
    .X(_14947_));
 sky130_fd_sc_hd__xnor2_2 _25038_ (.A(_14943_),
    .B(_14947_),
    .Y(_14948_));
 sky130_fd_sc_hd__buf_1 _25039_ (.A(_14948_),
    .X(_14949_));
 sky130_fd_sc_hd__nor2_2 _25040_ (.A(_11578_),
    .B(_14949_),
    .Y(_14950_));
 sky130_fd_sc_hd__xnor2_2 _25041_ (.A(_14939_),
    .B(_14950_),
    .Y(_14951_));
 sky130_fd_sc_hd__or4_2 _25042_ (.A(_12223_),
    .B(_12457_),
    .C(_14386_),
    .D(_13891_),
    .X(_14952_));
 sky130_fd_sc_hd__a22o_2 _25043_ (.A1(_12460_),
    .A2(_13542_),
    .B1(_13888_),
    .B2(_12225_),
    .X(_14954_));
 sky130_fd_sc_hd__nand2_2 _25044_ (.A(_14952_),
    .B(_14954_),
    .Y(_14955_));
 sky130_fd_sc_hd__nand2_2 _25045_ (.A(_14388_),
    .B(_14391_),
    .Y(_14956_));
 sky130_fd_sc_hd__xnor2_2 _25046_ (.A(_14955_),
    .B(_14956_),
    .Y(_14957_));
 sky130_fd_sc_hd__o21a_2 _25047_ (.A1(_14616_),
    .A2(_14617_),
    .B1(_14614_),
    .X(_14958_));
 sky130_fd_sc_hd__xnor2_2 _25048_ (.A(_14957_),
    .B(_14958_),
    .Y(_14959_));
 sky130_fd_sc_hd__xor2_2 _25049_ (.A(_14951_),
    .B(_14959_),
    .X(_14960_));
 sky130_fd_sc_hd__o21a_2 _25050_ (.A1(_14936_),
    .A2(_14937_),
    .B1(_14960_),
    .X(_14961_));
 sky130_fd_sc_hd__nor3_2 _25051_ (.A(_14936_),
    .B(_14937_),
    .C(_14960_),
    .Y(_14962_));
 sky130_fd_sc_hd__nor2_2 _25052_ (.A(_14961_),
    .B(_14962_),
    .Y(_14963_));
 sky130_fd_sc_hd__xnor2_2 _25053_ (.A(_14935_),
    .B(_14963_),
    .Y(_14965_));
 sky130_fd_sc_hd__or2_2 _25054_ (.A(_14639_),
    .B(_14642_),
    .X(_14966_));
 sky130_fd_sc_hd__o21ai_2 _25055_ (.A1(_14651_),
    .A2(_14653_),
    .B1(_14647_),
    .Y(_14967_));
 sky130_fd_sc_hd__nor2_2 _25056_ (.A(_12773_),
    .B(_13241_),
    .Y(_14968_));
 sky130_fd_sc_hd__xnor2_2 _25057_ (.A(_14632_),
    .B(_14968_),
    .Y(_14969_));
 sky130_fd_sc_hd__o21a_2 _25058_ (.A1(_14343_),
    .A2(_14625_),
    .B1(_14969_),
    .X(_14970_));
 sky130_fd_sc_hd__nor3_2 _25059_ (.A(_14343_),
    .B(_14625_),
    .C(_14969_),
    .Y(_14971_));
 sky130_fd_sc_hd__or2_2 _25060_ (.A(_14970_),
    .B(_14971_),
    .X(_14972_));
 sky130_fd_sc_hd__xor2_2 _25061_ (.A(_14967_),
    .B(_14972_),
    .X(_14973_));
 sky130_fd_sc_hd__a21oi_2 _25062_ (.A1(_14633_),
    .A2(_14966_),
    .B1(_14973_),
    .Y(_14974_));
 sky130_fd_sc_hd__and3_2 _25063_ (.A(_14633_),
    .B(_14966_),
    .C(_14973_),
    .X(_14976_));
 sky130_fd_sc_hd__nor2_2 _25064_ (.A(_14974_),
    .B(_14976_),
    .Y(_14977_));
 sky130_fd_sc_hd__buf_1 _25065_ (.A(_12248_),
    .X(_14978_));
 sky130_fd_sc_hd__or4_2 _25066_ (.A(_13926_),
    .B(_14978_),
    .C(_13842_),
    .D(_13934_),
    .X(_14979_));
 sky130_fd_sc_hd__buf_1 _25067_ (.A(_12242_),
    .X(_14980_));
 sky130_fd_sc_hd__a22o_2 _25068_ (.A1(_14980_),
    .A2(_13845_),
    .B1(_13938_),
    .B2(_14649_),
    .X(_14981_));
 sky130_fd_sc_hd__nand2_2 _25069_ (.A(_14979_),
    .B(_14981_),
    .Y(_14982_));
 sky130_fd_sc_hd__buf_1 _25070_ (.A(_13502_),
    .X(_14983_));
 sky130_fd_sc_hd__nor2_2 _25071_ (.A(_14356_),
    .B(_14983_),
    .Y(_14984_));
 sky130_fd_sc_hd__xnor2_2 _25072_ (.A(_14982_),
    .B(_14984_),
    .Y(_14985_));
 sky130_fd_sc_hd__nand2_2 _25073_ (.A(_14367_),
    .B(_14368_),
    .Y(_14987_));
 sky130_fd_sc_hd__buf_1 _25074_ (.A(_14987_),
    .X(_14988_));
 sky130_fd_sc_hd__nor2_2 _25075_ (.A(_11793_),
    .B(_14988_),
    .Y(_14989_));
 sky130_fd_sc_hd__a21o_2 _25076_ (.A1(iX[13]),
    .A2(iX[45]),
    .B1(_14660_),
    .X(_14990_));
 sky130_fd_sc_hd__nand2_2 _25077_ (.A(iX[14]),
    .B(iX[46]),
    .Y(_14991_));
 sky130_fd_sc_hd__or2_2 _25078_ (.A(iX[14]),
    .B(iX[46]),
    .X(_14992_));
 sky130_fd_sc_hd__nand2_2 _25079_ (.A(_14991_),
    .B(_14992_),
    .Y(_14993_));
 sky130_fd_sc_hd__o21bai_2 _25080_ (.A1(_14662_),
    .A2(_14990_),
    .B1_N(_14993_),
    .Y(_14994_));
 sky130_fd_sc_hd__buf_2 _25081_ (.A(_14994_),
    .X(_14995_));
 sky130_fd_sc_hd__or3b_4 _25082_ (.A(_14662_),
    .B(_14990_),
    .C_N(_14993_),
    .X(_14996_));
 sky130_fd_sc_hd__nand2_2 _25083_ (.A(_14995_),
    .B(_14996_),
    .Y(_14998_));
 sky130_fd_sc_hd__nor3_2 _25084_ (.A(_14659_),
    .B(_14660_),
    .C(_14662_),
    .Y(_14999_));
 sky130_fd_sc_hd__a32o_2 _25085_ (.A1(_11380_),
    .A2(_14995_),
    .A3(_14996_),
    .B1(_11585_),
    .B2(_14999_),
    .X(_15000_));
 sky130_fd_sc_hd__o31a_2 _25086_ (.A1(_11576_),
    .A2(_14663_),
    .A3(_14998_),
    .B1(_15000_),
    .X(_15001_));
 sky130_fd_sc_hd__xor2_2 _25087_ (.A(_14989_),
    .B(_15001_),
    .X(_15002_));
 sky130_fd_sc_hd__or3_2 _25088_ (.A(_14659_),
    .B(_14660_),
    .C(_14662_),
    .X(_15003_));
 sky130_fd_sc_hd__buf_1 _25089_ (.A(_15003_),
    .X(_15004_));
 sky130_fd_sc_hd__buf_1 _25090_ (.A(_15004_),
    .X(_15005_));
 sky130_fd_sc_hd__nor2_2 _25091_ (.A(_11567_),
    .B(_15005_),
    .Y(_15006_));
 sky130_fd_sc_hd__nor2_2 _25092_ (.A(_14655_),
    .B(_14664_),
    .Y(_15007_));
 sky130_fd_sc_hd__a21oi_2 _25093_ (.A1(_14369_),
    .A2(_15006_),
    .B1(_15007_),
    .Y(_15009_));
 sky130_fd_sc_hd__xnor2_2 _25094_ (.A(_15002_),
    .B(_15009_),
    .Y(_15010_));
 sky130_fd_sc_hd__xnor2_2 _25095_ (.A(_14985_),
    .B(_15010_),
    .Y(_15011_));
 sky130_fd_sc_hd__and2_2 _25096_ (.A(_14654_),
    .B(_14667_),
    .X(_15012_));
 sky130_fd_sc_hd__a21oi_2 _25097_ (.A1(_14665_),
    .A2(_14666_),
    .B1(_15012_),
    .Y(_15013_));
 sky130_fd_sc_hd__xor2_2 _25098_ (.A(_15011_),
    .B(_15013_),
    .X(_15014_));
 sky130_fd_sc_hd__xnor2_2 _25099_ (.A(_14977_),
    .B(_15014_),
    .Y(_15015_));
 sky130_fd_sc_hd__and2b_2 _25100_ (.A_N(_14669_),
    .B(_14671_),
    .X(_15016_));
 sky130_fd_sc_hd__a21oi_2 _25101_ (.A1(_14645_),
    .A2(_14672_),
    .B1(_15016_),
    .Y(_15017_));
 sky130_fd_sc_hd__xor2_2 _25102_ (.A(_15015_),
    .B(_15017_),
    .X(_15018_));
 sky130_fd_sc_hd__xnor2_2 _25103_ (.A(_14965_),
    .B(_15018_),
    .Y(_15020_));
 sky130_fd_sc_hd__and2b_2 _25104_ (.A_N(_14673_),
    .B(_14675_),
    .X(_15021_));
 sky130_fd_sc_hd__a21oi_2 _25105_ (.A1(_14623_),
    .A2(_14676_),
    .B1(_15021_),
    .Y(_15022_));
 sky130_fd_sc_hd__xnor2_2 _25106_ (.A(_15020_),
    .B(_15022_),
    .Y(_15023_));
 sky130_fd_sc_hd__xor2_2 _25107_ (.A(_14934_),
    .B(_15023_),
    .X(_15024_));
 sky130_fd_sc_hd__and2b_2 _25108_ (.A_N(_14681_),
    .B(_14683_),
    .X(_15025_));
 sky130_fd_sc_hd__o21ba_2 _25109_ (.A1(_14677_),
    .A2(_14680_),
    .B1_N(_15025_),
    .X(_15026_));
 sky130_fd_sc_hd__xnor2_2 _25110_ (.A(_15024_),
    .B(_15026_),
    .Y(_15027_));
 sky130_fd_sc_hd__xnor2_2 _25111_ (.A(_14927_),
    .B(_15027_),
    .Y(_15028_));
 sky130_fd_sc_hd__and3_2 _25112_ (.A(_14926_),
    .B(_14689_),
    .C(_15028_),
    .X(_15029_));
 sky130_fd_sc_hd__nor2_2 _25113_ (.A(_14689_),
    .B(_15028_),
    .Y(_15031_));
 sky130_fd_sc_hd__or2_2 _25114_ (.A(_14926_),
    .B(_15028_),
    .X(_15032_));
 sky130_fd_sc_hd__nor3b_2 _25115_ (.A(_15029_),
    .B(_15031_),
    .C_N(_15032_),
    .Y(_15033_));
 sky130_fd_sc_hd__nor2_2 _25116_ (.A(_14589_),
    .B(_14688_),
    .Y(_15034_));
 sky130_fd_sc_hd__a211o_2 _25117_ (.A1(_14425_),
    .A2(_14426_),
    .B1(_15034_),
    .C1(_14587_),
    .X(_15035_));
 sky130_fd_sc_hd__nand2_2 _25118_ (.A(_14692_),
    .B(_15035_),
    .Y(_15036_));
 sky130_fd_sc_hd__xor2_2 _25119_ (.A(_15033_),
    .B(_15036_),
    .X(_15037_));
 sky130_fd_sc_hd__a2bb2o_2 _25120_ (.A1_N(_14492_),
    .A2_N(_14583_),
    .B1(_14585_),
    .B2(_14513_),
    .X(_15038_));
 sky130_fd_sc_hd__nor2_2 _25121_ (.A(_14490_),
    .B(_14583_),
    .Y(_15039_));
 sky130_fd_sc_hd__and2b_2 _25122_ (.A_N(_14579_),
    .B(_14577_),
    .X(_15040_));
 sky130_fd_sc_hd__inv_2 _25123_ (.A(_15040_),
    .Y(_15042_));
 sky130_fd_sc_hd__nand2_2 _25124_ (.A(_14547_),
    .B(_14549_),
    .Y(_15043_));
 sky130_fd_sc_hd__or2b_2 _25125_ (.A(_14524_),
    .B_N(_14523_),
    .X(_15044_));
 sky130_fd_sc_hd__nand2_2 _25126_ (.A(_14525_),
    .B(_14531_),
    .Y(_15045_));
 sky130_fd_sc_hd__and4_2 _25127_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[43]),
    .D(iX[44]),
    .X(_15046_));
 sky130_fd_sc_hd__a22oi_2 _25128_ (.A1(iY[35]),
    .A2(iX[43]),
    .B1(iX[44]),
    .B2(iY[34]),
    .Y(_15047_));
 sky130_fd_sc_hd__nor2_2 _25129_ (.A(_15046_),
    .B(_15047_),
    .Y(_15048_));
 sky130_fd_sc_hd__nand2_2 _25130_ (.A(iY[33]),
    .B(iX[45]),
    .Y(_15049_));
 sky130_fd_sc_hd__xnor2_2 _25131_ (.A(_15048_),
    .B(_15049_),
    .Y(_15050_));
 sky130_fd_sc_hd__o21ba_2 _25132_ (.A1(_14520_),
    .A2(_14522_),
    .B1_N(_14519_),
    .X(_15051_));
 sky130_fd_sc_hd__xnor2_2 _25133_ (.A(_15050_),
    .B(_15051_),
    .Y(_15053_));
 sky130_fd_sc_hd__and4_2 _25134_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[42]),
    .D(iX[46]),
    .X(_15054_));
 sky130_fd_sc_hd__a22oi_2 _25135_ (.A1(iY[36]),
    .A2(iX[42]),
    .B1(iX[46]),
    .B2(iY[32]),
    .Y(_15055_));
 sky130_fd_sc_hd__nor2_2 _25136_ (.A(_15054_),
    .B(_15055_),
    .Y(_15056_));
 sky130_fd_sc_hd__nand2_2 _25137_ (.A(iY[37]),
    .B(iX[41]),
    .Y(_15057_));
 sky130_fd_sc_hd__xnor2_2 _25138_ (.A(_15056_),
    .B(_15057_),
    .Y(_15058_));
 sky130_fd_sc_hd__xnor2_2 _25139_ (.A(_15053_),
    .B(_15058_),
    .Y(_15059_));
 sky130_fd_sc_hd__a21o_2 _25140_ (.A1(_15044_),
    .A2(_15045_),
    .B1(_15059_),
    .X(_15060_));
 sky130_fd_sc_hd__nand3_2 _25141_ (.A(_15044_),
    .B(_15045_),
    .C(_15059_),
    .Y(_15061_));
 sky130_fd_sc_hd__o21ba_2 _25142_ (.A1(_14539_),
    .A2(_14541_),
    .B1_N(_14538_),
    .X(_15062_));
 sky130_fd_sc_hd__o21ba_2 _25143_ (.A1(_14528_),
    .A2(_14530_),
    .B1_N(_14527_),
    .X(_15064_));
 sky130_fd_sc_hd__and4_2 _25144_ (.A(iY[38]),
    .B(iX[39]),
    .C(iY[39]),
    .D(iX[40]),
    .X(_15065_));
 sky130_fd_sc_hd__a22oi_2 _25145_ (.A1(iX[39]),
    .A2(iY[39]),
    .B1(iX[40]),
    .B2(iY[38]),
    .Y(_15066_));
 sky130_fd_sc_hd__nor2_2 _25146_ (.A(_15065_),
    .B(_15066_),
    .Y(_15067_));
 sky130_fd_sc_hd__nand2_2 _25147_ (.A(iX[38]),
    .B(iY[40]),
    .Y(_15068_));
 sky130_fd_sc_hd__xnor2_2 _25148_ (.A(_15067_),
    .B(_15068_),
    .Y(_15069_));
 sky130_fd_sc_hd__xnor2_2 _25149_ (.A(_15064_),
    .B(_15069_),
    .Y(_15070_));
 sky130_fd_sc_hd__xnor2_2 _25150_ (.A(_15062_),
    .B(_15070_),
    .Y(_15071_));
 sky130_fd_sc_hd__nand3_2 _25151_ (.A(_15060_),
    .B(_15061_),
    .C(_15071_),
    .Y(_15072_));
 sky130_fd_sc_hd__a21o_2 _25152_ (.A1(_15060_),
    .A2(_15061_),
    .B1(_15071_),
    .X(_15073_));
 sky130_fd_sc_hd__nand2_2 _25153_ (.A(_15072_),
    .B(_15073_),
    .Y(_15075_));
 sky130_fd_sc_hd__a21o_2 _25154_ (.A1(_14533_),
    .A2(_14545_),
    .B1(_15075_),
    .X(_15076_));
 sky130_fd_sc_hd__nand3_2 _25155_ (.A(_14533_),
    .B(_14545_),
    .C(_15075_),
    .Y(_15077_));
 sky130_fd_sc_hd__or2b_2 _25156_ (.A(_14563_),
    .B_N(_14562_),
    .X(_15078_));
 sky130_fd_sc_hd__or2b_2 _25157_ (.A(_14556_),
    .B_N(_14564_),
    .X(_15079_));
 sky130_fd_sc_hd__or2b_2 _25158_ (.A(_14536_),
    .B_N(_14542_),
    .X(_15080_));
 sky130_fd_sc_hd__or2b_2 _25159_ (.A(_14535_),
    .B_N(_14543_),
    .X(_15081_));
 sky130_fd_sc_hd__and4_2 _25160_ (.A(iX[33]),
    .B(iX[34]),
    .C(iY[44]),
    .D(iY[45]),
    .X(_15082_));
 sky130_fd_sc_hd__a22oi_2 _25161_ (.A1(iX[34]),
    .A2(iY[44]),
    .B1(iY[45]),
    .B2(iX[33]),
    .Y(_15083_));
 sky130_fd_sc_hd__nor2_2 _25162_ (.A(_15082_),
    .B(_15083_),
    .Y(_15084_));
 sky130_fd_sc_hd__nand2_2 _25163_ (.A(iX[32]),
    .B(iY[46]),
    .Y(_15086_));
 sky130_fd_sc_hd__xnor2_2 _25164_ (.A(_15084_),
    .B(_15086_),
    .Y(_15087_));
 sky130_fd_sc_hd__and4_2 _25165_ (.A(iX[36]),
    .B(iX[37]),
    .C(iY[41]),
    .D(iY[42]),
    .X(_15088_));
 sky130_fd_sc_hd__a22oi_2 _25166_ (.A1(iX[37]),
    .A2(iY[41]),
    .B1(iY[42]),
    .B2(iX[36]),
    .Y(_15089_));
 sky130_fd_sc_hd__nor2_2 _25167_ (.A(_15088_),
    .B(_15089_),
    .Y(_15090_));
 sky130_fd_sc_hd__nand2_2 _25168_ (.A(iX[35]),
    .B(iY[43]),
    .Y(_15091_));
 sky130_fd_sc_hd__xnor2_2 _25169_ (.A(_15090_),
    .B(_15091_),
    .Y(_15092_));
 sky130_fd_sc_hd__o21ba_2 _25170_ (.A1(_14558_),
    .A2(_14561_),
    .B1_N(_14557_),
    .X(_15093_));
 sky130_fd_sc_hd__xnor2_2 _25171_ (.A(_15092_),
    .B(_15093_),
    .Y(_15094_));
 sky130_fd_sc_hd__and2_2 _25172_ (.A(_15087_),
    .B(_15094_),
    .X(_15095_));
 sky130_fd_sc_hd__nor2_2 _25173_ (.A(_15087_),
    .B(_15094_),
    .Y(_15097_));
 sky130_fd_sc_hd__or2_2 _25174_ (.A(_15095_),
    .B(_15097_),
    .X(_15098_));
 sky130_fd_sc_hd__a21o_2 _25175_ (.A1(_15080_),
    .A2(_15081_),
    .B1(_15098_),
    .X(_15099_));
 sky130_fd_sc_hd__inv_2 _25176_ (.A(_15099_),
    .Y(_15100_));
 sky130_fd_sc_hd__and3_2 _25177_ (.A(_15080_),
    .B(_15081_),
    .C(_15098_),
    .X(_15101_));
 sky130_fd_sc_hd__a211o_2 _25178_ (.A1(_15078_),
    .A2(_15079_),
    .B1(_15100_),
    .C1(_15101_),
    .X(_15102_));
 sky130_fd_sc_hd__o211ai_2 _25179_ (.A1(_15100_),
    .A2(_15101_),
    .B1(_15078_),
    .C1(_15079_),
    .Y(_15103_));
 sky130_fd_sc_hd__nand4_2 _25180_ (.A(_15076_),
    .B(_15077_),
    .C(_15102_),
    .D(_15103_),
    .Y(_15104_));
 sky130_fd_sc_hd__a22o_2 _25181_ (.A1(_15076_),
    .A2(_15077_),
    .B1(_15102_),
    .B2(_15103_),
    .X(_15105_));
 sky130_fd_sc_hd__nand2_2 _25182_ (.A(_15104_),
    .B(_15105_),
    .Y(_15106_));
 sky130_fd_sc_hd__a21o_2 _25183_ (.A1(_15043_),
    .A2(_14571_),
    .B1(_15106_),
    .X(_15108_));
 sky130_fd_sc_hd__nand3_2 _25184_ (.A(_15043_),
    .B(_14571_),
    .C(_15106_),
    .Y(_15109_));
 sky130_fd_sc_hd__o21ai_2 _25185_ (.A1(_14566_),
    .A2(_14568_),
    .B1(_14555_),
    .Y(_15110_));
 sky130_fd_sc_hd__or3_2 _25186_ (.A(_14555_),
    .B(_14566_),
    .C(_14568_),
    .X(_15111_));
 sky130_fd_sc_hd__and2_2 _25187_ (.A(_15110_),
    .B(_15111_),
    .X(_15112_));
 sky130_fd_sc_hd__a21o_2 _25188_ (.A1(_15108_),
    .A2(_15109_),
    .B1(_15112_),
    .X(_15113_));
 sky130_fd_sc_hd__nand3_2 _25189_ (.A(_15108_),
    .B(_15109_),
    .C(_15112_),
    .Y(_15114_));
 sky130_fd_sc_hd__nand2_2 _25190_ (.A(_15113_),
    .B(_15114_),
    .Y(_15115_));
 sky130_fd_sc_hd__o21ba_2 _25191_ (.A1(_14574_),
    .A2(_14576_),
    .B1_N(_14573_),
    .X(_15116_));
 sky130_fd_sc_hd__xnor2_2 _25192_ (.A(_15115_),
    .B(_15116_),
    .Y(_15117_));
 sky130_fd_sc_hd__xnor2_2 _25193_ (.A(_15042_),
    .B(_15117_),
    .Y(_15119_));
 sky130_fd_sc_hd__nand2_2 _25194_ (.A(_14581_),
    .B(_15119_),
    .Y(_15120_));
 sky130_fd_sc_hd__or3_2 _25195_ (.A(_14490_),
    .B(_14583_),
    .C(_15119_),
    .X(_15121_));
 sky130_fd_sc_hd__or2_2 _25196_ (.A(_14581_),
    .B(_15119_),
    .X(_15122_));
 sky130_fd_sc_hd__o211a_2 _25197_ (.A1(_15039_),
    .A2(_15120_),
    .B1(_15121_),
    .C1(_15122_),
    .X(_15123_));
 sky130_fd_sc_hd__xor2_2 _25198_ (.A(_15038_),
    .B(_15123_),
    .X(_15124_));
 sky130_fd_sc_hd__xor2_2 _25199_ (.A(_15037_),
    .B(_15124_),
    .X(_15125_));
 sky130_fd_sc_hd__xor2_2 _25200_ (.A(oO[14]),
    .B(_15125_),
    .X(_15126_));
 sky130_fd_sc_hd__and2b_2 _25201_ (.A_N(oO[13]),
    .B(_14695_),
    .X(_15127_));
 sky130_fd_sc_hd__a21oi_2 _25202_ (.A1(_14586_),
    .A2(_14694_),
    .B1(_15127_),
    .Y(_15128_));
 sky130_fd_sc_hd__xor2_2 _25203_ (.A(_15126_),
    .B(_15128_),
    .X(_15130_));
 sky130_fd_sc_hd__or2_2 _25204_ (.A(_14696_),
    .B(_14698_),
    .X(_15131_));
 sky130_fd_sc_hd__o21ai_2 _25205_ (.A1(_14699_),
    .A2(_14702_),
    .B1(_15131_),
    .Y(_15132_));
 sky130_fd_sc_hd__xor2_2 _25206_ (.A(_15130_),
    .B(_15132_),
    .X(_15133_));
 sky130_fd_sc_hd__xor2_2 _25207_ (.A(_14925_),
    .B(_15133_),
    .X(_15134_));
 sky130_fd_sc_hd__inv_2 _25208_ (.A(_15134_),
    .Y(_15135_));
 sky130_fd_sc_hd__inv_2 _25209_ (.A(_14816_),
    .Y(_15136_));
 sky130_fd_sc_hd__o21ai_2 _25210_ (.A1(_15136_),
    .A2(_14821_),
    .B1(_14818_),
    .Y(_15137_));
 sky130_fd_sc_hd__xnor2_2 _25211_ (.A(_15135_),
    .B(_15137_),
    .Y(oO[46]));
 sky130_fd_sc_hd__or2b_2 _25212_ (.A(_14925_),
    .B_N(_15133_),
    .X(_15138_));
 sky130_fd_sc_hd__o311ai_2 _25213_ (.A1(_14820_),
    .A2(_14510_),
    .A3(_15136_),
    .B1(_14818_),
    .C1(_15135_),
    .Y(_15140_));
 sky130_fd_sc_hd__or2_2 _25214_ (.A(_15037_),
    .B(_15124_),
    .X(_15141_));
 sky130_fd_sc_hd__or2b_2 _25215_ (.A(oO[14]),
    .B_N(_15125_),
    .X(_15142_));
 sky130_fd_sc_hd__a31o_4 _25216_ (.A1(_14692_),
    .A2(_15033_),
    .A3(_15035_),
    .B1(_15031_),
    .X(_15143_));
 sky130_fd_sc_hd__and2b_2 _25217_ (.A_N(_15026_),
    .B(_15024_),
    .X(_15144_));
 sky130_fd_sc_hd__a21o_2 _25218_ (.A1(_14935_),
    .A2(_14963_),
    .B1(_14961_),
    .X(_15145_));
 sky130_fd_sc_hd__or2_2 _25219_ (.A(_14609_),
    .B(_14938_),
    .X(_15146_));
 sky130_fd_sc_hd__a21boi_2 _25220_ (.A1(_14939_),
    .A2(_14950_),
    .B1_N(_15146_),
    .Y(_15147_));
 sky130_fd_sc_hd__nor2_2 _25221_ (.A(iY[15]),
    .B(iY[47]),
    .Y(_15148_));
 sky130_fd_sc_hd__nand2_2 _25222_ (.A(iY[15]),
    .B(iY[47]),
    .Y(_15149_));
 sky130_fd_sc_hd__nor2b_2 _25223_ (.A(_15148_),
    .B_N(_15149_),
    .Y(_15151_));
 sky130_fd_sc_hd__a21oi_2 _25224_ (.A1(_14943_),
    .A2(_14947_),
    .B1(_14940_),
    .Y(_15152_));
 sky130_fd_sc_hd__xor2_2 _25225_ (.A(_15151_),
    .B(_15152_),
    .X(_15153_));
 sky130_fd_sc_hd__buf_1 _25226_ (.A(_15153_),
    .X(_15154_));
 sky130_fd_sc_hd__buf_1 _25227_ (.A(_15154_),
    .X(_15155_));
 sky130_fd_sc_hd__or3_2 _25228_ (.A(_11579_),
    .B(_15147_),
    .C(_15155_),
    .X(_15156_));
 sky130_fd_sc_hd__o21ai_2 _25229_ (.A1(_11579_),
    .A2(_15155_),
    .B1(_15147_),
    .Y(_15157_));
 sky130_fd_sc_hd__and2_2 _25230_ (.A(_15156_),
    .B(_15157_),
    .X(_15158_));
 sky130_fd_sc_hd__xnor2_2 _25231_ (.A(_15145_),
    .B(_15158_),
    .Y(_15159_));
 sky130_fd_sc_hd__nor2_2 _25232_ (.A(_15015_),
    .B(_15017_),
    .Y(_15160_));
 sky130_fd_sc_hd__and2b_2 _25233_ (.A_N(_14965_),
    .B(_15018_),
    .X(_15162_));
 sky130_fd_sc_hd__or2_2 _25234_ (.A(_14957_),
    .B(_14958_),
    .X(_15163_));
 sky130_fd_sc_hd__or2_2 _25235_ (.A(_14951_),
    .B(_14959_),
    .X(_15164_));
 sky130_fd_sc_hd__and2b_2 _25236_ (.A_N(_14972_),
    .B(_14967_),
    .X(_15165_));
 sky130_fd_sc_hd__and3b_2 _25237_ (.A_N(_14938_),
    .B(_14605_),
    .C(_14388_),
    .X(_15166_));
 sky130_fd_sc_hd__buf_6 _25238_ (.A(_11827_),
    .X(_15167_));
 sky130_fd_sc_hd__nand2_2 _25239_ (.A(_14407_),
    .B(_14408_),
    .Y(_15168_));
 sky130_fd_sc_hd__or2_2 _25240_ (.A(_14601_),
    .B(_14603_),
    .X(_15169_));
 sky130_fd_sc_hd__o22a_2 _25241_ (.A1(_15167_),
    .A2(_15168_),
    .B1(_15169_),
    .B2(_12468_),
    .X(_15170_));
 sky130_fd_sc_hd__nor2_2 _25242_ (.A(_15166_),
    .B(_15170_),
    .Y(_15171_));
 sky130_fd_sc_hd__buf_1 _25243_ (.A(_14948_),
    .X(_15173_));
 sky130_fd_sc_hd__nor2_2 _25244_ (.A(_11570_),
    .B(_15173_),
    .Y(_15174_));
 sky130_fd_sc_hd__xnor2_2 _25245_ (.A(_15171_),
    .B(_15174_),
    .Y(_15175_));
 sky130_fd_sc_hd__or4_2 _25246_ (.A(_12457_),
    .B(_14343_),
    .C(_14386_),
    .D(_13891_),
    .X(_15176_));
 sky130_fd_sc_hd__a22o_2 _25247_ (.A1(_12816_),
    .A2(_13542_),
    .B1(_13887_),
    .B2(_12460_),
    .X(_15177_));
 sky130_fd_sc_hd__nand2_2 _25248_ (.A(_15176_),
    .B(_15177_),
    .Y(_15178_));
 sky130_fd_sc_hd__nand2_2 _25249_ (.A(_14628_),
    .B(_14391_),
    .Y(_15179_));
 sky130_fd_sc_hd__xnor2_2 _25250_ (.A(_15178_),
    .B(_15179_),
    .Y(_15180_));
 sky130_fd_sc_hd__o21a_2 _25251_ (.A1(_14955_),
    .A2(_14956_),
    .B1(_14952_),
    .X(_15181_));
 sky130_fd_sc_hd__xnor2_2 _25252_ (.A(_15180_),
    .B(_15181_),
    .Y(_15182_));
 sky130_fd_sc_hd__or2_2 _25253_ (.A(_15175_),
    .B(_15182_),
    .X(_15184_));
 sky130_fd_sc_hd__nand2_2 _25254_ (.A(_15175_),
    .B(_15182_),
    .Y(_15185_));
 sky130_fd_sc_hd__and2_2 _25255_ (.A(_15184_),
    .B(_15185_),
    .X(_15186_));
 sky130_fd_sc_hd__o21a_2 _25256_ (.A1(_15165_),
    .A2(_14974_),
    .B1(_15186_),
    .X(_15187_));
 sky130_fd_sc_hd__nor3_2 _25257_ (.A(_15165_),
    .B(_14974_),
    .C(_15186_),
    .Y(_15188_));
 sky130_fd_sc_hd__a211oi_2 _25258_ (.A1(_15163_),
    .A2(_15164_),
    .B1(_15187_),
    .C1(_15188_),
    .Y(_15189_));
 sky130_fd_sc_hd__o211a_2 _25259_ (.A1(_15187_),
    .A2(_15188_),
    .B1(_15163_),
    .C1(_15164_),
    .X(_15190_));
 sky130_fd_sc_hd__or2_2 _25260_ (.A(_15011_),
    .B(_15013_),
    .X(_15191_));
 sky130_fd_sc_hd__nand2_2 _25261_ (.A(_14977_),
    .B(_15014_),
    .Y(_15192_));
 sky130_fd_sc_hd__a21o_2 _25262_ (.A1(_14632_),
    .A2(_14968_),
    .B1(_14971_),
    .X(_15193_));
 sky130_fd_sc_hd__a21bo_2 _25263_ (.A1(_14981_),
    .A2(_14984_),
    .B1_N(_14979_),
    .X(_15195_));
 sky130_fd_sc_hd__or3b_2 _25264_ (.A(_12850_),
    .B(_13502_),
    .C_N(_14968_),
    .X(_15196_));
 sky130_fd_sc_hd__a22o_2 _25265_ (.A1(_12846_),
    .A2(_13244_),
    .B1(_13496_),
    .B2(_14634_),
    .X(_15197_));
 sky130_fd_sc_hd__nand2_2 _25266_ (.A(_15196_),
    .B(_15197_),
    .Y(_15198_));
 sky130_fd_sc_hd__nor2_2 _25267_ (.A(_14357_),
    .B(_14641_),
    .Y(_15199_));
 sky130_fd_sc_hd__xnor2_2 _25268_ (.A(_15198_),
    .B(_15199_),
    .Y(_15200_));
 sky130_fd_sc_hd__nand2_2 _25269_ (.A(_15195_),
    .B(_15200_),
    .Y(_15201_));
 sky130_fd_sc_hd__or2_2 _25270_ (.A(_15195_),
    .B(_15200_),
    .X(_15202_));
 sky130_fd_sc_hd__and2_2 _25271_ (.A(_15201_),
    .B(_15202_),
    .X(_15203_));
 sky130_fd_sc_hd__xnor2_2 _25272_ (.A(_15193_),
    .B(_15203_),
    .Y(_15204_));
 sky130_fd_sc_hd__or4_2 _25273_ (.A(_13926_),
    .B(_12248_),
    .C(_13934_),
    .D(_14987_),
    .X(_15206_));
 sky130_fd_sc_hd__and2_2 _25274_ (.A(_14367_),
    .B(_14368_),
    .X(_15207_));
 sky130_fd_sc_hd__buf_1 _25275_ (.A(_15207_),
    .X(_15208_));
 sky130_fd_sc_hd__a22o_2 _25276_ (.A1(_14980_),
    .A2(_13938_),
    .B1(_15208_),
    .B2(_14649_),
    .X(_15209_));
 sky130_fd_sc_hd__nand2_2 _25277_ (.A(_15206_),
    .B(_15209_),
    .Y(_15210_));
 sky130_fd_sc_hd__buf_1 _25278_ (.A(_13842_),
    .X(_15211_));
 sky130_fd_sc_hd__nor2_2 _25279_ (.A(_14356_),
    .B(_15211_),
    .Y(_15212_));
 sky130_fd_sc_hd__xnor2_2 _25280_ (.A(_15210_),
    .B(_15212_),
    .Y(_15213_));
 sky130_fd_sc_hd__nor2_2 _25281_ (.A(_11793_),
    .B(_15005_),
    .Y(_15214_));
 sky130_fd_sc_hd__nor2_2 _25282_ (.A(iX[15]),
    .B(iX[47]),
    .Y(_15215_));
 sky130_fd_sc_hd__nand2_2 _25283_ (.A(iX[15]),
    .B(iX[47]),
    .Y(_15217_));
 sky130_fd_sc_hd__or2b_2 _25284_ (.A(_15215_),
    .B_N(_15217_),
    .X(_15218_));
 sky130_fd_sc_hd__and3_2 _25285_ (.A(_14991_),
    .B(_14995_),
    .C(_15218_),
    .X(_15219_));
 sky130_fd_sc_hd__a21oi_2 _25286_ (.A1(_14991_),
    .A2(_14995_),
    .B1(_15218_),
    .Y(_15220_));
 sky130_fd_sc_hd__and3_2 _25287_ (.A(_11583_),
    .B(_14995_),
    .C(_14996_),
    .X(_15221_));
 sky130_fd_sc_hd__or4b_4 _25288_ (.A(_11566_),
    .B(_15219_),
    .C(_15220_),
    .D_N(_15221_),
    .X(_15222_));
 sky130_fd_sc_hd__nand3_2 _25289_ (.A(_14991_),
    .B(_14995_),
    .C(_15218_),
    .Y(_15223_));
 sky130_fd_sc_hd__buf_1 _25290_ (.A(_15223_),
    .X(_15224_));
 sky130_fd_sc_hd__a21o_2 _25291_ (.A1(_14991_),
    .A2(_14995_),
    .B1(_15218_),
    .X(_15225_));
 sky130_fd_sc_hd__buf_2 _25292_ (.A(_15225_),
    .X(_15226_));
 sky130_fd_sc_hd__a31o_2 _25293_ (.A1(_11381_),
    .A2(_15224_),
    .A3(_15226_),
    .B1(_15221_),
    .X(_15228_));
 sky130_fd_sc_hd__nand3_2 _25294_ (.A(_15214_),
    .B(_15222_),
    .C(_15228_),
    .Y(_15229_));
 sky130_fd_sc_hd__a21o_2 _25295_ (.A1(_15222_),
    .A2(_15228_),
    .B1(_15214_),
    .X(_15230_));
 sky130_fd_sc_hd__a22o_2 _25296_ (.A1(_15006_),
    .A2(_15221_),
    .B1(_15001_),
    .B2(_14989_),
    .X(_15231_));
 sky130_fd_sc_hd__nand3_2 _25297_ (.A(_15229_),
    .B(_15230_),
    .C(_15231_),
    .Y(_15232_));
 sky130_fd_sc_hd__a21o_2 _25298_ (.A1(_15229_),
    .A2(_15230_),
    .B1(_15231_),
    .X(_15233_));
 sky130_fd_sc_hd__nand3_2 _25299_ (.A(_15213_),
    .B(_15232_),
    .C(_15233_),
    .Y(_15234_));
 sky130_fd_sc_hd__a21o_2 _25300_ (.A1(_15232_),
    .A2(_15233_),
    .B1(_15213_),
    .X(_15235_));
 sky130_fd_sc_hd__and2b_2 _25301_ (.A_N(_15009_),
    .B(_15002_),
    .X(_15236_));
 sky130_fd_sc_hd__a21o_2 _25302_ (.A1(_14985_),
    .A2(_15010_),
    .B1(_15236_),
    .X(_15237_));
 sky130_fd_sc_hd__and3_2 _25303_ (.A(_15234_),
    .B(_15235_),
    .C(_15237_),
    .X(_15239_));
 sky130_fd_sc_hd__a21oi_2 _25304_ (.A1(_15234_),
    .A2(_15235_),
    .B1(_15237_),
    .Y(_15240_));
 sky130_fd_sc_hd__nor3_2 _25305_ (.A(_15204_),
    .B(_15239_),
    .C(_15240_),
    .Y(_15241_));
 sky130_fd_sc_hd__o21a_2 _25306_ (.A1(_15239_),
    .A2(_15240_),
    .B1(_15204_),
    .X(_15242_));
 sky130_fd_sc_hd__a211oi_2 _25307_ (.A1(_15191_),
    .A2(_15192_),
    .B1(_15241_),
    .C1(_15242_),
    .Y(_15243_));
 sky130_fd_sc_hd__o211a_2 _25308_ (.A1(_15241_),
    .A2(_15242_),
    .B1(_15191_),
    .C1(_15192_),
    .X(_15244_));
 sky130_fd_sc_hd__or4_4 _25309_ (.A(_15189_),
    .B(_15190_),
    .C(_15243_),
    .D(_15244_),
    .X(_15245_));
 sky130_fd_sc_hd__o22ai_2 _25310_ (.A1(_15189_),
    .A2(_15190_),
    .B1(_15243_),
    .B2(_15244_),
    .Y(_15246_));
 sky130_fd_sc_hd__o211a_2 _25311_ (.A1(_15160_),
    .A2(_15162_),
    .B1(_15245_),
    .C1(_15246_),
    .X(_15247_));
 sky130_fd_sc_hd__a211oi_2 _25312_ (.A1(_15245_),
    .A2(_15246_),
    .B1(_15160_),
    .C1(_15162_),
    .Y(_15248_));
 sky130_fd_sc_hd__or3_2 _25313_ (.A(_15159_),
    .B(_15247_),
    .C(_15248_),
    .X(_15250_));
 sky130_fd_sc_hd__o21ai_2 _25314_ (.A1(_15247_),
    .A2(_15248_),
    .B1(_15159_),
    .Y(_15251_));
 sky130_fd_sc_hd__and2b_2 _25315_ (.A_N(_15022_),
    .B(_15020_),
    .X(_15252_));
 sky130_fd_sc_hd__a21o_2 _25316_ (.A1(_14934_),
    .A2(_15023_),
    .B1(_15252_),
    .X(_15253_));
 sky130_fd_sc_hd__nand3_2 _25317_ (.A(_15250_),
    .B(_15251_),
    .C(_15253_),
    .Y(_15254_));
 sky130_fd_sc_hd__a21o_2 _25318_ (.A1(_15250_),
    .A2(_15251_),
    .B1(_15253_),
    .X(_15255_));
 sky130_fd_sc_hd__nand3_2 _25319_ (.A(_14932_),
    .B(_15254_),
    .C(_15255_),
    .Y(_15256_));
 sky130_fd_sc_hd__a21o_2 _25320_ (.A1(_15254_),
    .A2(_15255_),
    .B1(_14932_),
    .X(_15257_));
 sky130_fd_sc_hd__and3_2 _25321_ (.A(_15144_),
    .B(_15256_),
    .C(_15257_),
    .X(_15258_));
 sky130_fd_sc_hd__a21o_2 _25322_ (.A1(_15256_),
    .A2(_15257_),
    .B1(_15144_),
    .X(_15259_));
 sky130_fd_sc_hd__or2b_2 _25323_ (.A(_15258_),
    .B_N(_15259_),
    .X(_15261_));
 sky130_fd_sc_hd__and2_2 _25324_ (.A(_14927_),
    .B(_15027_),
    .X(_15262_));
 sky130_fd_sc_hd__or2b_2 _25325_ (.A(_15262_),
    .B_N(_15032_),
    .X(_15263_));
 sky130_fd_sc_hd__xnor2_2 _25326_ (.A(_15261_),
    .B(_15263_),
    .Y(_15264_));
 sky130_fd_sc_hd__xnor2_2 _25327_ (.A(_15143_),
    .B(_15264_),
    .Y(_15265_));
 sky130_fd_sc_hd__a21bo_2 _25328_ (.A1(_15038_),
    .A2(_15123_),
    .B1_N(_15121_),
    .X(_15266_));
 sky130_fd_sc_hd__or2_2 _25329_ (.A(_15115_),
    .B(_15116_),
    .X(_15267_));
 sky130_fd_sc_hd__or2b_2 _25330_ (.A(_15051_),
    .B_N(_15050_),
    .X(_15268_));
 sky130_fd_sc_hd__nand2_2 _25331_ (.A(_15053_),
    .B(_15058_),
    .Y(_15269_));
 sky130_fd_sc_hd__and4_2 _25332_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[44]),
    .D(iX[45]),
    .X(_15270_));
 sky130_fd_sc_hd__a22oi_2 _25333_ (.A1(iY[35]),
    .A2(iX[44]),
    .B1(iX[45]),
    .B2(iY[34]),
    .Y(_15272_));
 sky130_fd_sc_hd__nor2_2 _25334_ (.A(_15270_),
    .B(_15272_),
    .Y(_15273_));
 sky130_fd_sc_hd__nand2_2 _25335_ (.A(iY[33]),
    .B(iX[46]),
    .Y(_15274_));
 sky130_fd_sc_hd__xnor2_2 _25336_ (.A(_15273_),
    .B(_15274_),
    .Y(_15275_));
 sky130_fd_sc_hd__o21ba_2 _25337_ (.A1(_15047_),
    .A2(_15049_),
    .B1_N(_15046_),
    .X(_15276_));
 sky130_fd_sc_hd__xnor2_2 _25338_ (.A(_15275_),
    .B(_15276_),
    .Y(_15277_));
 sky130_fd_sc_hd__and4_2 _25339_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[43]),
    .D(iX[47]),
    .X(_15278_));
 sky130_fd_sc_hd__a22oi_2 _25340_ (.A1(iY[36]),
    .A2(iX[43]),
    .B1(iX[47]),
    .B2(iY[32]),
    .Y(_15279_));
 sky130_fd_sc_hd__nor2_2 _25341_ (.A(_15278_),
    .B(_15279_),
    .Y(_15280_));
 sky130_fd_sc_hd__nand2_2 _25342_ (.A(iY[37]),
    .B(iX[42]),
    .Y(_15281_));
 sky130_fd_sc_hd__xnor2_2 _25343_ (.A(_15280_),
    .B(_15281_),
    .Y(_15283_));
 sky130_fd_sc_hd__xnor2_2 _25344_ (.A(_15277_),
    .B(_15283_),
    .Y(_15284_));
 sky130_fd_sc_hd__a21o_2 _25345_ (.A1(_15268_),
    .A2(_15269_),
    .B1(_15284_),
    .X(_15285_));
 sky130_fd_sc_hd__nand3_2 _25346_ (.A(_15268_),
    .B(_15269_),
    .C(_15284_),
    .Y(_15286_));
 sky130_fd_sc_hd__o21ba_2 _25347_ (.A1(_15066_),
    .A2(_15068_),
    .B1_N(_15065_),
    .X(_15287_));
 sky130_fd_sc_hd__o21ba_2 _25348_ (.A1(_15055_),
    .A2(_15057_),
    .B1_N(_15054_),
    .X(_15288_));
 sky130_fd_sc_hd__and4_2 _25349_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[40]),
    .D(iX[41]),
    .X(_15289_));
 sky130_fd_sc_hd__a22oi_2 _25350_ (.A1(iY[39]),
    .A2(iX[40]),
    .B1(iX[41]),
    .B2(iY[38]),
    .Y(_15290_));
 sky130_fd_sc_hd__nor2_2 _25351_ (.A(_15289_),
    .B(_15290_),
    .Y(_15291_));
 sky130_fd_sc_hd__nand2_2 _25352_ (.A(iX[39]),
    .B(iY[40]),
    .Y(_15292_));
 sky130_fd_sc_hd__xnor2_2 _25353_ (.A(_15291_),
    .B(_15292_),
    .Y(_15294_));
 sky130_fd_sc_hd__xnor2_2 _25354_ (.A(_15288_),
    .B(_15294_),
    .Y(_15295_));
 sky130_fd_sc_hd__xnor2_2 _25355_ (.A(_15287_),
    .B(_15295_),
    .Y(_15296_));
 sky130_fd_sc_hd__nand3_2 _25356_ (.A(_15285_),
    .B(_15286_),
    .C(_15296_),
    .Y(_15297_));
 sky130_fd_sc_hd__a21o_2 _25357_ (.A1(_15285_),
    .A2(_15286_),
    .B1(_15296_),
    .X(_15298_));
 sky130_fd_sc_hd__nand2_2 _25358_ (.A(_15297_),
    .B(_15298_),
    .Y(_15299_));
 sky130_fd_sc_hd__a21o_2 _25359_ (.A1(_15060_),
    .A2(_15072_),
    .B1(_15299_),
    .X(_15300_));
 sky130_fd_sc_hd__nand3_2 _25360_ (.A(_15060_),
    .B(_15072_),
    .C(_15299_),
    .Y(_15301_));
 sky130_fd_sc_hd__nand2_2 _25361_ (.A(_15300_),
    .B(_15301_),
    .Y(_15302_));
 sky130_fd_sc_hd__and2b_2 _25362_ (.A_N(_15093_),
    .B(_15092_),
    .X(_15303_));
 sky130_fd_sc_hd__or2b_2 _25363_ (.A(_15064_),
    .B_N(_15069_),
    .X(_15305_));
 sky130_fd_sc_hd__or2b_2 _25364_ (.A(_15062_),
    .B_N(_15070_),
    .X(_15306_));
 sky130_fd_sc_hd__and4_2 _25365_ (.A(iX[34]),
    .B(iX[35]),
    .C(iY[44]),
    .D(iY[45]),
    .X(_15307_));
 sky130_fd_sc_hd__a22oi_2 _25366_ (.A1(iX[35]),
    .A2(iY[44]),
    .B1(iY[45]),
    .B2(iX[34]),
    .Y(_15308_));
 sky130_fd_sc_hd__nor2_2 _25367_ (.A(_15307_),
    .B(_15308_),
    .Y(_15309_));
 sky130_fd_sc_hd__nand2_2 _25368_ (.A(iX[33]),
    .B(iY[46]),
    .Y(_15310_));
 sky130_fd_sc_hd__xnor2_2 _25369_ (.A(_15309_),
    .B(_15310_),
    .Y(_15311_));
 sky130_fd_sc_hd__and4_2 _25370_ (.A(iX[37]),
    .B(iX[38]),
    .C(iY[41]),
    .D(iY[42]),
    .X(_15312_));
 sky130_fd_sc_hd__a22oi_2 _25371_ (.A1(iX[38]),
    .A2(iY[41]),
    .B1(iY[42]),
    .B2(iX[37]),
    .Y(_15313_));
 sky130_fd_sc_hd__nor2_2 _25372_ (.A(_15312_),
    .B(_15313_),
    .Y(_15314_));
 sky130_fd_sc_hd__nand2_2 _25373_ (.A(iX[36]),
    .B(iY[43]),
    .Y(_15316_));
 sky130_fd_sc_hd__xnor2_2 _25374_ (.A(_15314_),
    .B(_15316_),
    .Y(_15317_));
 sky130_fd_sc_hd__o21ba_2 _25375_ (.A1(_15089_),
    .A2(_15091_),
    .B1_N(_15088_),
    .X(_15318_));
 sky130_fd_sc_hd__xnor2_2 _25376_ (.A(_15317_),
    .B(_15318_),
    .Y(_15319_));
 sky130_fd_sc_hd__and2_2 _25377_ (.A(_15311_),
    .B(_15319_),
    .X(_15320_));
 sky130_fd_sc_hd__nor2_2 _25378_ (.A(_15311_),
    .B(_15319_),
    .Y(_15321_));
 sky130_fd_sc_hd__or2_2 _25379_ (.A(_15320_),
    .B(_15321_),
    .X(_15322_));
 sky130_fd_sc_hd__a21o_2 _25380_ (.A1(_15305_),
    .A2(_15306_),
    .B1(_15322_),
    .X(_15323_));
 sky130_fd_sc_hd__nand3_2 _25381_ (.A(_15305_),
    .B(_15306_),
    .C(_15322_),
    .Y(_15324_));
 sky130_fd_sc_hd__o211ai_2 _25382_ (.A1(_15303_),
    .A2(_15095_),
    .B1(_15323_),
    .C1(_15324_),
    .Y(_15325_));
 sky130_fd_sc_hd__a211o_2 _25383_ (.A1(_15323_),
    .A2(_15324_),
    .B1(_15303_),
    .C1(_15095_),
    .X(_15327_));
 sky130_fd_sc_hd__nand2_2 _25384_ (.A(_15325_),
    .B(_15327_),
    .Y(_15328_));
 sky130_fd_sc_hd__xnor2_2 _25385_ (.A(_15302_),
    .B(_15328_),
    .Y(_15329_));
 sky130_fd_sc_hd__nand2_2 _25386_ (.A(_15076_),
    .B(_15104_),
    .Y(_15330_));
 sky130_fd_sc_hd__xor2_2 _25387_ (.A(_15329_),
    .B(_15330_),
    .X(_15331_));
 sky130_fd_sc_hd__o21ba_2 _25388_ (.A1(_15083_),
    .A2(_15086_),
    .B1_N(_15082_),
    .X(_15332_));
 sky130_fd_sc_hd__nand2_2 _25389_ (.A(iX[32]),
    .B(iY[47]),
    .Y(_15333_));
 sky130_fd_sc_hd__xnor2_2 _25390_ (.A(_15332_),
    .B(_15333_),
    .Y(_15334_));
 sky130_fd_sc_hd__a21o_2 _25391_ (.A1(_15099_),
    .A2(_15102_),
    .B1(_15334_),
    .X(_15335_));
 sky130_fd_sc_hd__nand3_2 _25392_ (.A(_15099_),
    .B(_15102_),
    .C(_15334_),
    .Y(_15336_));
 sky130_fd_sc_hd__and2_2 _25393_ (.A(_15335_),
    .B(_15336_),
    .X(_15338_));
 sky130_fd_sc_hd__xnor2_2 _25394_ (.A(_15331_),
    .B(_15338_),
    .Y(_15339_));
 sky130_fd_sc_hd__inv_2 _25395_ (.A(_15339_),
    .Y(_15340_));
 sky130_fd_sc_hd__a21oi_2 _25396_ (.A1(_15108_),
    .A2(_15114_),
    .B1(_15340_),
    .Y(_15341_));
 sky130_fd_sc_hd__and3_2 _25397_ (.A(_15108_),
    .B(_15114_),
    .C(_15340_),
    .X(_15342_));
 sky130_fd_sc_hd__nor3_2 _25398_ (.A(_15110_),
    .B(_15341_),
    .C(_15342_),
    .Y(_15343_));
 sky130_fd_sc_hd__o21a_2 _25399_ (.A1(_15341_),
    .A2(_15342_),
    .B1(_15110_),
    .X(_15344_));
 sky130_fd_sc_hd__or2_2 _25400_ (.A(_15343_),
    .B(_15344_),
    .X(_15345_));
 sky130_fd_sc_hd__xor2_2 _25401_ (.A(_15267_),
    .B(_15345_),
    .X(_15346_));
 sky130_fd_sc_hd__nor2_2 _25402_ (.A(_15042_),
    .B(_15117_),
    .Y(_15347_));
 sky130_fd_sc_hd__and2b_2 _25403_ (.A_N(_15347_),
    .B(_15122_),
    .X(_15349_));
 sky130_fd_sc_hd__xnor2_2 _25404_ (.A(_15346_),
    .B(_15349_),
    .Y(_15350_));
 sky130_fd_sc_hd__xor2_2 _25405_ (.A(_15266_),
    .B(_15350_),
    .X(_15351_));
 sky130_fd_sc_hd__xnor2_2 _25406_ (.A(_15265_),
    .B(_15351_),
    .Y(_15352_));
 sky130_fd_sc_hd__xnor2_2 _25407_ (.A(oO[15]),
    .B(_15352_),
    .Y(_15353_));
 sky130_fd_sc_hd__a21oi_2 _25408_ (.A1(_15141_),
    .A2(_15142_),
    .B1(_15353_),
    .Y(_15354_));
 sky130_fd_sc_hd__and3_2 _25409_ (.A(_15141_),
    .B(_15142_),
    .C(_15353_),
    .X(_15355_));
 sky130_fd_sc_hd__nor2_2 _25410_ (.A(_15354_),
    .B(_15355_),
    .Y(_15356_));
 sky130_fd_sc_hd__nor2_2 _25411_ (.A(_15126_),
    .B(_15128_),
    .Y(_15357_));
 sky130_fd_sc_hd__a21o_2 _25412_ (.A1(_15130_),
    .A2(_15132_),
    .B1(_15357_),
    .X(_15358_));
 sky130_fd_sc_hd__xnor2_2 _25413_ (.A(_15356_),
    .B(_15358_),
    .Y(_15360_));
 sky130_fd_sc_hd__o21a_2 _25414_ (.A1(_14799_),
    .A2(_14802_),
    .B1(_14912_),
    .X(_15361_));
 sky130_fd_sc_hd__and2b_2 _25415_ (.A_N(_14910_),
    .B(_14911_),
    .X(_15362_));
 sky130_fd_sc_hd__and2b_2 _25416_ (.A_N(_14830_),
    .B(_14829_),
    .X(_15363_));
 sky130_fd_sc_hd__nand2_2 _25417_ (.A(iY[16]),
    .B(iX[30]),
    .Y(_15364_));
 sky130_fd_sc_hd__nand2_2 _25418_ (.A(iY[17]),
    .B(iX[31]),
    .Y(_15365_));
 sky130_fd_sc_hd__a22o_2 _25419_ (.A1(iY[17]),
    .A2(iX[30]),
    .B1(iX[31]),
    .B2(iY[16]),
    .X(_15366_));
 sky130_fd_sc_hd__o21a_2 _25420_ (.A1(_15364_),
    .A2(_15365_),
    .B1(_15366_),
    .X(_15367_));
 sky130_fd_sc_hd__a31o_2 _25421_ (.A1(iY[17]),
    .A2(iX[29]),
    .A3(_14826_),
    .B1(_14825_),
    .X(_15368_));
 sky130_fd_sc_hd__nand2_2 _25422_ (.A(_15367_),
    .B(_15368_),
    .Y(_15369_));
 sky130_fd_sc_hd__or2_2 _25423_ (.A(_15367_),
    .B(_15368_),
    .X(_15371_));
 sky130_fd_sc_hd__and2_2 _25424_ (.A(_15369_),
    .B(_15371_),
    .X(_15372_));
 sky130_fd_sc_hd__nand2_2 _25425_ (.A(_15363_),
    .B(_15372_),
    .Y(_15373_));
 sky130_fd_sc_hd__or2_2 _25426_ (.A(_15363_),
    .B(_15372_),
    .X(_15374_));
 sky130_fd_sc_hd__nand2_2 _25427_ (.A(_15373_),
    .B(_15374_),
    .Y(_15375_));
 sky130_fd_sc_hd__and4_2 _25428_ (.A(iY[21]),
    .B(iY[22]),
    .C(iX[25]),
    .D(iX[26]),
    .X(_15376_));
 sky130_fd_sc_hd__a22oi_2 _25429_ (.A1(iY[22]),
    .A2(iX[25]),
    .B1(iX[26]),
    .B2(iY[21]),
    .Y(_15377_));
 sky130_fd_sc_hd__nor2_2 _25430_ (.A(_15376_),
    .B(_15377_),
    .Y(_15378_));
 sky130_fd_sc_hd__nand2_2 _25431_ (.A(iY[23]),
    .B(iX[24]),
    .Y(_15379_));
 sky130_fd_sc_hd__xnor2_2 _25432_ (.A(_15378_),
    .B(_15379_),
    .Y(_15380_));
 sky130_fd_sc_hd__and4_2 _25433_ (.A(iY[18]),
    .B(iY[19]),
    .C(iX[28]),
    .D(iX[29]),
    .X(_15381_));
 sky130_fd_sc_hd__a22oi_2 _25434_ (.A1(iY[19]),
    .A2(iX[28]),
    .B1(iX[29]),
    .B2(iY[18]),
    .Y(_15382_));
 sky130_fd_sc_hd__nor2_2 _25435_ (.A(_15381_),
    .B(_15382_),
    .Y(_15383_));
 sky130_fd_sc_hd__nand2_2 _25436_ (.A(iY[20]),
    .B(iX[27]),
    .Y(_15384_));
 sky130_fd_sc_hd__xnor2_2 _25437_ (.A(_15383_),
    .B(_15384_),
    .Y(_15385_));
 sky130_fd_sc_hd__o21ba_2 _25438_ (.A1(_14842_),
    .A2(_14845_),
    .B1_N(_14841_),
    .X(_15386_));
 sky130_fd_sc_hd__xnor2_2 _25439_ (.A(_15385_),
    .B(_15386_),
    .Y(_15387_));
 sky130_fd_sc_hd__and2_2 _25440_ (.A(_15380_),
    .B(_15387_),
    .X(_15388_));
 sky130_fd_sc_hd__nor2_2 _25441_ (.A(_15380_),
    .B(_15387_),
    .Y(_15389_));
 sky130_fd_sc_hd__or2_2 _25442_ (.A(_15388_),
    .B(_15389_),
    .X(_15390_));
 sky130_fd_sc_hd__or2_2 _25443_ (.A(_15375_),
    .B(_15390_),
    .X(_15392_));
 sky130_fd_sc_hd__nand2_2 _25444_ (.A(_15375_),
    .B(_15390_),
    .Y(_15393_));
 sky130_fd_sc_hd__nand2_2 _25445_ (.A(_15392_),
    .B(_15393_),
    .Y(_15394_));
 sky130_fd_sc_hd__a21oi_2 _25446_ (.A1(_14835_),
    .A2(_14852_),
    .B1(_14833_),
    .Y(_15395_));
 sky130_fd_sc_hd__xnor2_2 _25447_ (.A(_15394_),
    .B(_15395_),
    .Y(_15396_));
 sky130_fd_sc_hd__or2b_2 _25448_ (.A(_14866_),
    .B_N(_14864_),
    .X(_15397_));
 sky130_fd_sc_hd__and4_2 _25449_ (.A(iX[19]),
    .B(iX[20]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_15398_));
 sky130_fd_sc_hd__a22oi_2 _25450_ (.A1(iX[20]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[19]),
    .Y(_15399_));
 sky130_fd_sc_hd__nor2_2 _25451_ (.A(_15398_),
    .B(_15399_),
    .Y(_15400_));
 sky130_fd_sc_hd__nand2_2 _25452_ (.A(iX[18]),
    .B(iY[29]),
    .Y(_15401_));
 sky130_fd_sc_hd__xnor2_2 _25453_ (.A(_15400_),
    .B(_15401_),
    .Y(_15403_));
 sky130_fd_sc_hd__o21ba_2 _25454_ (.A1(_14861_),
    .A2(_14863_),
    .B1_N(_14860_),
    .X(_15404_));
 sky130_fd_sc_hd__xnor2_2 _25455_ (.A(_15403_),
    .B(_15404_),
    .Y(_15405_));
 sky130_fd_sc_hd__nand3_2 _25456_ (.A(iX[17]),
    .B(iY[30]),
    .C(_15405_),
    .Y(_15406_));
 sky130_fd_sc_hd__a21o_2 _25457_ (.A1(iX[17]),
    .A2(iY[30]),
    .B1(_15405_),
    .X(_15407_));
 sky130_fd_sc_hd__nand2_2 _25458_ (.A(_15406_),
    .B(_15407_),
    .Y(_15408_));
 sky130_fd_sc_hd__a21oi_2 _25459_ (.A1(_15397_),
    .A2(_14870_),
    .B1(_15408_),
    .Y(_15409_));
 sky130_fd_sc_hd__and3_2 _25460_ (.A(_15397_),
    .B(_14870_),
    .C(_15408_),
    .X(_15410_));
 sky130_fd_sc_hd__nor2_2 _25461_ (.A(_15409_),
    .B(_15410_),
    .Y(_15411_));
 sky130_fd_sc_hd__nand2_2 _25462_ (.A(iX[16]),
    .B(iY[31]),
    .Y(_15412_));
 sky130_fd_sc_hd__xnor2_2 _25463_ (.A(_15411_),
    .B(_15412_),
    .Y(_15414_));
 sky130_fd_sc_hd__or2b_2 _25464_ (.A(_14882_),
    .B_N(_14888_),
    .X(_15415_));
 sky130_fd_sc_hd__or2b_2 _25465_ (.A(_14881_),
    .B_N(_14889_),
    .X(_15416_));
 sky130_fd_sc_hd__and2b_2 _25466_ (.A_N(_14847_),
    .B(_14846_),
    .X(_15417_));
 sky130_fd_sc_hd__o21ba_2 _25467_ (.A1(_14884_),
    .A2(_14886_),
    .B1_N(_14883_),
    .X(_15418_));
 sky130_fd_sc_hd__o21ba_2 _25468_ (.A1(_14837_),
    .A2(_14839_),
    .B1_N(_14836_),
    .X(_15419_));
 sky130_fd_sc_hd__and4_2 _25469_ (.A(iX[22]),
    .B(iX[23]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_15420_));
 sky130_fd_sc_hd__a22oi_2 _25470_ (.A1(iX[23]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[22]),
    .Y(_15421_));
 sky130_fd_sc_hd__nor2_2 _25471_ (.A(_15420_),
    .B(_15421_),
    .Y(_15422_));
 sky130_fd_sc_hd__nand2_2 _25472_ (.A(iX[21]),
    .B(iY[26]),
    .Y(_15423_));
 sky130_fd_sc_hd__xnor2_2 _25473_ (.A(_15422_),
    .B(_15423_),
    .Y(_15425_));
 sky130_fd_sc_hd__xnor2_2 _25474_ (.A(_15419_),
    .B(_15425_),
    .Y(_15426_));
 sky130_fd_sc_hd__xnor2_2 _25475_ (.A(_15418_),
    .B(_15426_),
    .Y(_15427_));
 sky130_fd_sc_hd__o21a_2 _25476_ (.A1(_15417_),
    .A2(_14849_),
    .B1(_15427_),
    .X(_15428_));
 sky130_fd_sc_hd__nor3_2 _25477_ (.A(_15417_),
    .B(_14849_),
    .C(_15427_),
    .Y(_15429_));
 sky130_fd_sc_hd__a211oi_2 _25478_ (.A1(_15415_),
    .A2(_15416_),
    .B1(_15428_),
    .C1(_15429_),
    .Y(_15430_));
 sky130_fd_sc_hd__o211a_2 _25479_ (.A1(_15428_),
    .A2(_15429_),
    .B1(_15415_),
    .C1(_15416_),
    .X(_15431_));
 sky130_fd_sc_hd__nor2_2 _25480_ (.A(_14891_),
    .B(_14893_),
    .Y(_15432_));
 sky130_fd_sc_hd__or3_2 _25481_ (.A(_15430_),
    .B(_15431_),
    .C(_15432_),
    .X(_15433_));
 sky130_fd_sc_hd__o21ai_2 _25482_ (.A1(_15430_),
    .A2(_15431_),
    .B1(_15432_),
    .Y(_15434_));
 sky130_fd_sc_hd__nand3_2 _25483_ (.A(_15414_),
    .B(_15433_),
    .C(_15434_),
    .Y(_15436_));
 sky130_fd_sc_hd__a21o_2 _25484_ (.A1(_15433_),
    .A2(_15434_),
    .B1(_15414_),
    .X(_15437_));
 sky130_fd_sc_hd__and3_2 _25485_ (.A(_14855_),
    .B(_15436_),
    .C(_15437_),
    .X(_15438_));
 sky130_fd_sc_hd__a21oi_2 _25486_ (.A1(_15436_),
    .A2(_15437_),
    .B1(_14855_),
    .Y(_15439_));
 sky130_fd_sc_hd__a211oi_2 _25487_ (.A1(_14896_),
    .A2(_14899_),
    .B1(_15438_),
    .C1(_15439_),
    .Y(_15440_));
 sky130_fd_sc_hd__o211a_2 _25488_ (.A1(_15438_),
    .A2(_15439_),
    .B1(_14896_),
    .C1(_14899_),
    .X(_15441_));
 sky130_fd_sc_hd__or3_2 _25489_ (.A(_15396_),
    .B(_15440_),
    .C(_15441_),
    .X(_15442_));
 sky130_fd_sc_hd__o21ai_2 _25490_ (.A1(_15440_),
    .A2(_15441_),
    .B1(_15396_),
    .Y(_15443_));
 sky130_fd_sc_hd__o21ai_2 _25491_ (.A1(_14824_),
    .A2(_14857_),
    .B1(_14905_),
    .Y(_15444_));
 sky130_fd_sc_hd__nand3_2 _25492_ (.A(_15442_),
    .B(_15443_),
    .C(_15444_),
    .Y(_15445_));
 sky130_fd_sc_hd__a21o_2 _25493_ (.A1(_15442_),
    .A2(_15443_),
    .B1(_15444_),
    .X(_15447_));
 sky130_fd_sc_hd__o211ai_2 _25494_ (.A1(_14901_),
    .A2(_14903_),
    .B1(_15445_),
    .C1(_15447_),
    .Y(_15448_));
 sky130_fd_sc_hd__a211o_2 _25495_ (.A1(_15445_),
    .A2(_15447_),
    .B1(_14901_),
    .C1(_14903_),
    .X(_15449_));
 sky130_fd_sc_hd__o211a_2 _25496_ (.A1(_14907_),
    .A2(_15362_),
    .B1(_15448_),
    .C1(_15449_),
    .X(_15450_));
 sky130_fd_sc_hd__a211oi_2 _25497_ (.A1(_15448_),
    .A2(_15449_),
    .B1(_14907_),
    .C1(_15362_),
    .Y(_15451_));
 sky130_fd_sc_hd__nor2_2 _25498_ (.A(_15450_),
    .B(_15451_),
    .Y(_15452_));
 sky130_fd_sc_hd__a31o_2 _25499_ (.A1(iX[15]),
    .A2(iY[31]),
    .A3(_14874_),
    .B1(_14872_),
    .X(_15453_));
 sky130_fd_sc_hd__xor2_2 _25500_ (.A(_15452_),
    .B(_15453_),
    .X(_15454_));
 sky130_fd_sc_hd__or3_2 _25501_ (.A(_15361_),
    .B(_14915_),
    .C(_15454_),
    .X(_15455_));
 sky130_fd_sc_hd__o21ai_2 _25502_ (.A1(_15361_),
    .A2(_14915_),
    .B1(_15454_),
    .Y(_15456_));
 sky130_fd_sc_hd__nand2_2 _25503_ (.A(_15455_),
    .B(_15456_),
    .Y(_15458_));
 sky130_fd_sc_hd__a21oi_2 _25504_ (.A1(_14922_),
    .A2(_14924_),
    .B1(_14919_),
    .Y(_15459_));
 sky130_fd_sc_hd__xnor2_2 _25505_ (.A(_15458_),
    .B(_15459_),
    .Y(_15460_));
 sky130_fd_sc_hd__or2_2 _25506_ (.A(_15360_),
    .B(_15460_),
    .X(_15461_));
 sky130_fd_sc_hd__nand2_2 _25507_ (.A(_15360_),
    .B(_15460_),
    .Y(_15462_));
 sky130_fd_sc_hd__nand2_2 _25508_ (.A(_15461_),
    .B(_15462_),
    .Y(_15463_));
 sky130_fd_sc_hd__a21oi_2 _25509_ (.A1(_15138_),
    .A2(_15140_),
    .B1(_15463_),
    .Y(_15464_));
 sky130_fd_sc_hd__and3_2 _25510_ (.A(_15138_),
    .B(_15140_),
    .C(_15463_),
    .X(_15465_));
 sky130_fd_sc_hd__nor2_2 _25511_ (.A(_15464_),
    .B(_15465_),
    .Y(oO[47]));
 sky130_fd_sc_hd__a21o_2 _25512_ (.A1(_15138_),
    .A2(_15140_),
    .B1(_15463_),
    .X(_15466_));
 sky130_fd_sc_hd__and2_2 _25513_ (.A(_15461_),
    .B(_15466_),
    .X(_15468_));
 sky130_fd_sc_hd__inv_2 _25514_ (.A(_15458_),
    .Y(_15469_));
 sky130_fd_sc_hd__and4b_2 _25515_ (.A_N(_14328_),
    .B(_14813_),
    .C(_14922_),
    .D(_15469_),
    .X(_15470_));
 sky130_fd_sc_hd__nor4b_2 _25516_ (.A(_13220_),
    .B(_13483_),
    .C(_14331_),
    .D_N(_15470_),
    .Y(_15471_));
 sky130_fd_sc_hd__or2b_2 _25517_ (.A(_14332_),
    .B_N(_15470_),
    .X(_15472_));
 sky130_fd_sc_hd__a21bo_2 _25518_ (.A1(_13228_),
    .A2(_15471_),
    .B1_N(_15472_),
    .X(_15473_));
 sky130_fd_sc_hd__nand2_2 _25519_ (.A(_14922_),
    .B(_15469_),
    .Y(_15474_));
 sky130_fd_sc_hd__nand2_2 _25520_ (.A(_14919_),
    .B(_15455_),
    .Y(_15475_));
 sky130_fd_sc_hd__o211ai_2 _25521_ (.A1(_14923_),
    .A2(_15474_),
    .B1(_15475_),
    .C1(_15456_),
    .Y(_15476_));
 sky130_fd_sc_hd__or2_2 _25522_ (.A(_15473_),
    .B(_15476_),
    .X(_15477_));
 sky130_fd_sc_hd__o21ba_2 _25523_ (.A1(_15410_),
    .A2(_15412_),
    .B1_N(_15409_),
    .X(_15479_));
 sky130_fd_sc_hd__nor2_2 _25524_ (.A(_14708_),
    .B(_15365_),
    .Y(_15480_));
 sky130_fd_sc_hd__xor2_2 _25525_ (.A(_15369_),
    .B(_15480_),
    .X(_15481_));
 sky130_fd_sc_hd__and4_2 _25526_ (.A(iY[21]),
    .B(iY[22]),
    .C(iX[26]),
    .D(iX[27]),
    .X(_15482_));
 sky130_fd_sc_hd__a22oi_2 _25527_ (.A1(iY[22]),
    .A2(iX[26]),
    .B1(iX[27]),
    .B2(iY[21]),
    .Y(_15483_));
 sky130_fd_sc_hd__nor2_2 _25528_ (.A(_15482_),
    .B(_15483_),
    .Y(_15484_));
 sky130_fd_sc_hd__nand2_2 _25529_ (.A(iY[23]),
    .B(iX[25]),
    .Y(_15485_));
 sky130_fd_sc_hd__xnor2_2 _25530_ (.A(_15484_),
    .B(_15485_),
    .Y(_15486_));
 sky130_fd_sc_hd__and2_2 _25531_ (.A(iY[19]),
    .B(iX[30]),
    .X(_15487_));
 sky130_fd_sc_hd__and3_2 _25532_ (.A(iY[18]),
    .B(iX[29]),
    .C(_15487_),
    .X(_15488_));
 sky130_fd_sc_hd__a22oi_2 _25533_ (.A1(iY[19]),
    .A2(iX[29]),
    .B1(iX[30]),
    .B2(iY[18]),
    .Y(_15490_));
 sky130_fd_sc_hd__nor2_2 _25534_ (.A(_15488_),
    .B(_15490_),
    .Y(_15491_));
 sky130_fd_sc_hd__nand2_2 _25535_ (.A(iY[20]),
    .B(iX[28]),
    .Y(_15492_));
 sky130_fd_sc_hd__xnor2_2 _25536_ (.A(_15491_),
    .B(_15492_),
    .Y(_15493_));
 sky130_fd_sc_hd__o21ba_2 _25537_ (.A1(_15382_),
    .A2(_15384_),
    .B1_N(_15381_),
    .X(_15494_));
 sky130_fd_sc_hd__xnor2_2 _25538_ (.A(_15493_),
    .B(_15494_),
    .Y(_15495_));
 sky130_fd_sc_hd__and2_2 _25539_ (.A(_15486_),
    .B(_15495_),
    .X(_15496_));
 sky130_fd_sc_hd__nor2_2 _25540_ (.A(_15486_),
    .B(_15495_),
    .Y(_15497_));
 sky130_fd_sc_hd__or2_2 _25541_ (.A(_15496_),
    .B(_15497_),
    .X(_15498_));
 sky130_fd_sc_hd__nor2_2 _25542_ (.A(_15481_),
    .B(_15498_),
    .Y(_15499_));
 sky130_fd_sc_hd__and2_2 _25543_ (.A(_15481_),
    .B(_15498_),
    .X(_15501_));
 sky130_fd_sc_hd__a211o_2 _25544_ (.A1(_15373_),
    .A2(_15392_),
    .B1(_15499_),
    .C1(_15501_),
    .X(_15502_));
 sky130_fd_sc_hd__o211ai_2 _25545_ (.A1(_15499_),
    .A2(_15501_),
    .B1(_15373_),
    .C1(_15392_),
    .Y(_15503_));
 sky130_fd_sc_hd__or2_2 _25546_ (.A(_15394_),
    .B(_15395_),
    .X(_15504_));
 sky130_fd_sc_hd__or2b_2 _25547_ (.A(_15404_),
    .B_N(_15403_),
    .X(_15505_));
 sky130_fd_sc_hd__and4_2 _25548_ (.A(iX[20]),
    .B(iX[21]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_15506_));
 sky130_fd_sc_hd__a22oi_2 _25549_ (.A1(iX[21]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[20]),
    .Y(_15507_));
 sky130_fd_sc_hd__nor2_2 _25550_ (.A(_15506_),
    .B(_15507_),
    .Y(_15508_));
 sky130_fd_sc_hd__nand2_2 _25551_ (.A(iX[19]),
    .B(iY[29]),
    .Y(_15509_));
 sky130_fd_sc_hd__xnor2_2 _25552_ (.A(_15508_),
    .B(_15509_),
    .Y(_15510_));
 sky130_fd_sc_hd__o21ba_2 _25553_ (.A1(_15399_),
    .A2(_15401_),
    .B1_N(_15398_),
    .X(_15512_));
 sky130_fd_sc_hd__xnor2_2 _25554_ (.A(_15510_),
    .B(_15512_),
    .Y(_15513_));
 sky130_fd_sc_hd__nand3_2 _25555_ (.A(iX[18]),
    .B(iY[30]),
    .C(_15513_),
    .Y(_15514_));
 sky130_fd_sc_hd__a21o_2 _25556_ (.A1(iX[18]),
    .A2(iY[30]),
    .B1(_15513_),
    .X(_15515_));
 sky130_fd_sc_hd__nand2_2 _25557_ (.A(_15514_),
    .B(_15515_),
    .Y(_15516_));
 sky130_fd_sc_hd__a21o_2 _25558_ (.A1(_15505_),
    .A2(_15406_),
    .B1(_15516_),
    .X(_15517_));
 sky130_fd_sc_hd__nand3_2 _25559_ (.A(_15505_),
    .B(_15406_),
    .C(_15516_),
    .Y(_15518_));
 sky130_fd_sc_hd__nand2_2 _25560_ (.A(_15517_),
    .B(_15518_),
    .Y(_15519_));
 sky130_fd_sc_hd__nand2_2 _25561_ (.A(iX[17]),
    .B(iY[31]),
    .Y(_15520_));
 sky130_fd_sc_hd__nand2_2 _25562_ (.A(_15519_),
    .B(_15520_),
    .Y(_15521_));
 sky130_fd_sc_hd__or2_2 _25563_ (.A(_15519_),
    .B(_15520_),
    .X(_15523_));
 sky130_fd_sc_hd__and2_2 _25564_ (.A(_15521_),
    .B(_15523_),
    .X(_15524_));
 sky130_fd_sc_hd__or2b_2 _25565_ (.A(_15419_),
    .B_N(_15425_),
    .X(_15525_));
 sky130_fd_sc_hd__or2b_2 _25566_ (.A(_15418_),
    .B_N(_15426_),
    .X(_15526_));
 sky130_fd_sc_hd__and2b_2 _25567_ (.A_N(_15386_),
    .B(_15385_),
    .X(_15527_));
 sky130_fd_sc_hd__o21ba_2 _25568_ (.A1(_15421_),
    .A2(_15423_),
    .B1_N(_15420_),
    .X(_15528_));
 sky130_fd_sc_hd__o21ba_2 _25569_ (.A1(_15377_),
    .A2(_15379_),
    .B1_N(_15376_),
    .X(_15529_));
 sky130_fd_sc_hd__and4_2 _25570_ (.A(iX[23]),
    .B(iX[24]),
    .C(iY[24]),
    .D(iY[25]),
    .X(_15530_));
 sky130_fd_sc_hd__a22oi_2 _25571_ (.A1(iX[24]),
    .A2(iY[24]),
    .B1(iY[25]),
    .B2(iX[23]),
    .Y(_15531_));
 sky130_fd_sc_hd__nor2_2 _25572_ (.A(_15530_),
    .B(_15531_),
    .Y(_15532_));
 sky130_fd_sc_hd__nand2_2 _25573_ (.A(iX[22]),
    .B(iY[26]),
    .Y(_15534_));
 sky130_fd_sc_hd__xnor2_2 _25574_ (.A(_15532_),
    .B(_15534_),
    .Y(_15535_));
 sky130_fd_sc_hd__xnor2_2 _25575_ (.A(_15529_),
    .B(_15535_),
    .Y(_15536_));
 sky130_fd_sc_hd__xnor2_2 _25576_ (.A(_15528_),
    .B(_15536_),
    .Y(_15537_));
 sky130_fd_sc_hd__o21a_2 _25577_ (.A1(_15527_),
    .A2(_15388_),
    .B1(_15537_),
    .X(_15538_));
 sky130_fd_sc_hd__nor3_2 _25578_ (.A(_15527_),
    .B(_15388_),
    .C(_15537_),
    .Y(_15539_));
 sky130_fd_sc_hd__a211oi_2 _25579_ (.A1(_15525_),
    .A2(_15526_),
    .B1(_15538_),
    .C1(_15539_),
    .Y(_15540_));
 sky130_fd_sc_hd__o211a_2 _25580_ (.A1(_15538_),
    .A2(_15539_),
    .B1(_15525_),
    .C1(_15526_),
    .X(_15541_));
 sky130_fd_sc_hd__nor2_2 _25581_ (.A(_15428_),
    .B(_15430_),
    .Y(_15542_));
 sky130_fd_sc_hd__or3_2 _25582_ (.A(_15540_),
    .B(_15541_),
    .C(_15542_),
    .X(_15543_));
 sky130_fd_sc_hd__o21ai_2 _25583_ (.A1(_15540_),
    .A2(_15541_),
    .B1(_15542_),
    .Y(_15545_));
 sky130_fd_sc_hd__and3_2 _25584_ (.A(_15524_),
    .B(_15543_),
    .C(_15545_),
    .X(_15546_));
 sky130_fd_sc_hd__a21oi_2 _25585_ (.A1(_15543_),
    .A2(_15545_),
    .B1(_15524_),
    .Y(_15547_));
 sky130_fd_sc_hd__or3_2 _25586_ (.A(_15504_),
    .B(_15546_),
    .C(_15547_),
    .X(_15548_));
 sky130_fd_sc_hd__o21ai_2 _25587_ (.A1(_15546_),
    .A2(_15547_),
    .B1(_15504_),
    .Y(_15549_));
 sky130_fd_sc_hd__nand2_2 _25588_ (.A(_15548_),
    .B(_15549_),
    .Y(_15550_));
 sky130_fd_sc_hd__a21o_2 _25589_ (.A1(_15433_),
    .A2(_15436_),
    .B1(_15550_),
    .X(_15551_));
 sky130_fd_sc_hd__nand3_2 _25590_ (.A(_15433_),
    .B(_15436_),
    .C(_15550_),
    .Y(_15552_));
 sky130_fd_sc_hd__and4_2 _25591_ (.A(_15502_),
    .B(_15503_),
    .C(_15551_),
    .D(_15552_),
    .X(_15553_));
 sky130_fd_sc_hd__a22oi_2 _25592_ (.A1(_15502_),
    .A2(_15503_),
    .B1(_15551_),
    .B2(_15552_),
    .Y(_15554_));
 sky130_fd_sc_hd__or3_2 _25593_ (.A(_15442_),
    .B(_15553_),
    .C(_15554_),
    .X(_15556_));
 sky130_fd_sc_hd__o21ai_2 _25594_ (.A1(_15553_),
    .A2(_15554_),
    .B1(_15442_),
    .Y(_15557_));
 sky130_fd_sc_hd__o211ai_2 _25595_ (.A1(_15438_),
    .A2(_15440_),
    .B1(_15556_),
    .C1(_15557_),
    .Y(_15558_));
 sky130_fd_sc_hd__a211o_2 _25596_ (.A1(_15556_),
    .A2(_15557_),
    .B1(_15438_),
    .C1(_15440_),
    .X(_15559_));
 sky130_fd_sc_hd__and2_2 _25597_ (.A(_15558_),
    .B(_15559_),
    .X(_15560_));
 sky130_fd_sc_hd__nand2_2 _25598_ (.A(_15445_),
    .B(_15448_),
    .Y(_15561_));
 sky130_fd_sc_hd__nand2_2 _25599_ (.A(_15560_),
    .B(_15561_),
    .Y(_15562_));
 sky130_fd_sc_hd__or2_2 _25600_ (.A(_15560_),
    .B(_15561_),
    .X(_15563_));
 sky130_fd_sc_hd__and2_2 _25601_ (.A(_15562_),
    .B(_15563_),
    .X(_15564_));
 sky130_fd_sc_hd__or2b_2 _25602_ (.A(_15479_),
    .B_N(_15564_),
    .X(_15565_));
 sky130_fd_sc_hd__or2b_2 _25603_ (.A(_15564_),
    .B_N(_15479_),
    .X(_15567_));
 sky130_fd_sc_hd__nand2_2 _25604_ (.A(_15565_),
    .B(_15567_),
    .Y(_15568_));
 sky130_fd_sc_hd__a21oi_2 _25605_ (.A1(_15452_),
    .A2(_15453_),
    .B1(_15450_),
    .Y(_15569_));
 sky130_fd_sc_hd__nor2_2 _25606_ (.A(_15568_),
    .B(_15569_),
    .Y(_15570_));
 sky130_fd_sc_hd__and2_2 _25607_ (.A(_15568_),
    .B(_15569_),
    .X(_15571_));
 sky130_fd_sc_hd__nor2_2 _25608_ (.A(_15570_),
    .B(_15571_),
    .Y(_15572_));
 sky130_fd_sc_hd__nand2_2 _25609_ (.A(_15477_),
    .B(_15572_),
    .Y(_15573_));
 sky130_fd_sc_hd__or2_2 _25610_ (.A(_15477_),
    .B(_15572_),
    .X(_15574_));
 sky130_fd_sc_hd__and2_2 _25611_ (.A(_15573_),
    .B(_15574_),
    .X(_15575_));
 sky130_fd_sc_hd__or2_2 _25612_ (.A(_15265_),
    .B(_15351_),
    .X(_15576_));
 sky130_fd_sc_hd__o21a_2 _25613_ (.A1(oO[15]),
    .A2(_15352_),
    .B1(_15576_),
    .X(_15578_));
 sky130_fd_sc_hd__a2bb2o_2 _25614_ (.A1_N(_15032_),
    .A2_N(_15261_),
    .B1(_15264_),
    .B2(_15143_),
    .X(_15579_));
 sky130_fd_sc_hd__a21bo_2 _25615_ (.A1(_14932_),
    .A2(_15255_),
    .B1_N(_15254_),
    .X(_15580_));
 sky130_fd_sc_hd__and2_2 _25616_ (.A(_15145_),
    .B(_15158_),
    .X(_15581_));
 sky130_fd_sc_hd__nor3_2 _25617_ (.A(_15159_),
    .B(_15247_),
    .C(_15248_),
    .Y(_15582_));
 sky130_fd_sc_hd__and2_2 _25618_ (.A(_15171_),
    .B(_15174_),
    .X(_15583_));
 sky130_fd_sc_hd__or2_2 _25619_ (.A(_15166_),
    .B(_15583_),
    .X(_15584_));
 sky130_fd_sc_hd__xnor2_2 _25620_ (.A(_15151_),
    .B(_15152_),
    .Y(_15585_));
 sky130_fd_sc_hd__buf_1 _25621_ (.A(_15585_),
    .X(_15586_));
 sky130_fd_sc_hd__and3_2 _25622_ (.A(_14943_),
    .B(_14944_),
    .C(_15151_),
    .X(_15587_));
 sky130_fd_sc_hd__nand2_2 _25623_ (.A(iY[14]),
    .B(iY[46]),
    .Y(_15589_));
 sky130_fd_sc_hd__a21oi_2 _25624_ (.A1(_15589_),
    .A2(_15149_),
    .B1(_15148_),
    .Y(_15590_));
 sky130_fd_sc_hd__a31o_2 _25625_ (.A1(_14943_),
    .A2(_14946_),
    .A3(_15151_),
    .B1(_15590_),
    .X(_15591_));
 sky130_fd_sc_hd__a21o_2 _25626_ (.A1(_14402_),
    .A2(_15587_),
    .B1(_15591_),
    .X(_15592_));
 sky130_fd_sc_hd__and2_2 _25627_ (.A(iY[16]),
    .B(iY[48]),
    .X(_15593_));
 sky130_fd_sc_hd__nor2_2 _25628_ (.A(iY[16]),
    .B(iY[48]),
    .Y(_15594_));
 sky130_fd_sc_hd__nor2_2 _25629_ (.A(_15593_),
    .B(_15594_),
    .Y(_15595_));
 sky130_fd_sc_hd__xnor2_2 _25630_ (.A(_15592_),
    .B(_15595_),
    .Y(_15596_));
 sky130_fd_sc_hd__buf_1 _25631_ (.A(_15596_),
    .X(_15597_));
 sky130_fd_sc_hd__buf_1 _25632_ (.A(_15597_),
    .X(_15598_));
 sky130_fd_sc_hd__nor2_2 _25633_ (.A(_11570_),
    .B(_15598_),
    .Y(_15600_));
 sky130_fd_sc_hd__and3_2 _25634_ (.A(_11374_),
    .B(_15586_),
    .C(_15600_),
    .X(_15601_));
 sky130_fd_sc_hd__o22a_2 _25635_ (.A1(_11571_),
    .A2(_15155_),
    .B1(_15598_),
    .B2(_11578_),
    .X(_15602_));
 sky130_fd_sc_hd__or2_2 _25636_ (.A(_15601_),
    .B(_15602_),
    .X(_15603_));
 sky130_fd_sc_hd__xnor2_2 _25637_ (.A(_15584_),
    .B(_15603_),
    .Y(_15604_));
 sky130_fd_sc_hd__xnor2_2 _25638_ (.A(_15156_),
    .B(_15604_),
    .Y(_15605_));
 sky130_fd_sc_hd__o21a_2 _25639_ (.A1(_15187_),
    .A2(_15189_),
    .B1(_15605_),
    .X(_15606_));
 sky130_fd_sc_hd__nor3_2 _25640_ (.A(_15187_),
    .B(_15189_),
    .C(_15605_),
    .Y(_15607_));
 sky130_fd_sc_hd__nor2_2 _25641_ (.A(_15606_),
    .B(_15607_),
    .Y(_15608_));
 sky130_fd_sc_hd__a211o_2 _25642_ (.A1(_15191_),
    .A2(_15192_),
    .B1(_15241_),
    .C1(_15242_),
    .X(_15609_));
 sky130_fd_sc_hd__or2_2 _25643_ (.A(_15180_),
    .B(_15181_),
    .X(_15611_));
 sky130_fd_sc_hd__a21bo_2 _25644_ (.A1(_15193_),
    .A2(_15202_),
    .B1_N(_15201_),
    .X(_15612_));
 sky130_fd_sc_hd__nand2_2 _25645_ (.A(_14388_),
    .B(_14608_),
    .Y(_15613_));
 sky130_fd_sc_hd__nand2_2 _25646_ (.A(_14628_),
    .B(_14410_),
    .Y(_15614_));
 sky130_fd_sc_hd__xnor2_2 _25647_ (.A(_15613_),
    .B(_15614_),
    .Y(_15615_));
 sky130_fd_sc_hd__buf_1 _25648_ (.A(_12827_),
    .X(_15616_));
 sky130_fd_sc_hd__xor2_2 _25649_ (.A(_14943_),
    .B(_14947_),
    .X(_15617_));
 sky130_fd_sc_hd__nand2_2 _25650_ (.A(_15616_),
    .B(_15617_),
    .Y(_15618_));
 sky130_fd_sc_hd__xnor2_2 _25651_ (.A(_15615_),
    .B(_15618_),
    .Y(_15619_));
 sky130_fd_sc_hd__or4_2 _25652_ (.A(_14343_),
    .B(_12808_),
    .C(_14386_),
    .D(_13891_),
    .X(_15620_));
 sky130_fd_sc_hd__a22o_2 _25653_ (.A1(_13501_),
    .A2(_13543_),
    .B1(_13888_),
    .B2(_12816_),
    .X(_15622_));
 sky130_fd_sc_hd__nand2_2 _25654_ (.A(_15620_),
    .B(_15622_),
    .Y(_15623_));
 sky130_fd_sc_hd__buf_6 _25655_ (.A(_12460_),
    .X(_15624_));
 sky130_fd_sc_hd__nand2_2 _25656_ (.A(_15624_),
    .B(_14392_),
    .Y(_15625_));
 sky130_fd_sc_hd__xnor2_2 _25657_ (.A(_15623_),
    .B(_15625_),
    .Y(_15626_));
 sky130_fd_sc_hd__o21a_2 _25658_ (.A1(_15178_),
    .A2(_15179_),
    .B1(_15176_),
    .X(_15627_));
 sky130_fd_sc_hd__xnor2_2 _25659_ (.A(_15626_),
    .B(_15627_),
    .Y(_15628_));
 sky130_fd_sc_hd__xor2_2 _25660_ (.A(_15619_),
    .B(_15628_),
    .X(_15629_));
 sky130_fd_sc_hd__xnor2_2 _25661_ (.A(_15612_),
    .B(_15629_),
    .Y(_15630_));
 sky130_fd_sc_hd__a21oi_2 _25662_ (.A1(_15611_),
    .A2(_15184_),
    .B1(_15630_),
    .Y(_15631_));
 sky130_fd_sc_hd__and3_2 _25663_ (.A(_15611_),
    .B(_15184_),
    .C(_15630_),
    .X(_15633_));
 sky130_fd_sc_hd__nor2_2 _25664_ (.A(_15631_),
    .B(_15633_),
    .Y(_15634_));
 sky130_fd_sc_hd__a21bo_2 _25665_ (.A1(_15197_),
    .A2(_15199_),
    .B1_N(_15196_),
    .X(_15635_));
 sky130_fd_sc_hd__a21bo_2 _25666_ (.A1(_15209_),
    .A2(_15212_),
    .B1_N(_15206_),
    .X(_15636_));
 sky130_fd_sc_hd__nor2_2 _25667_ (.A(_12772_),
    .B(_13842_),
    .Y(_15637_));
 sky130_fd_sc_hd__and3_2 _25668_ (.A(_12846_),
    .B(_13496_),
    .C(_15637_),
    .X(_15638_));
 sky130_fd_sc_hd__a21oi_2 _25669_ (.A1(_12846_),
    .A2(_14648_),
    .B1(_15637_),
    .Y(_15639_));
 sky130_fd_sc_hd__nor2_2 _25670_ (.A(_15638_),
    .B(_15639_),
    .Y(_15640_));
 sky130_fd_sc_hd__nor2_2 _25671_ (.A(_14352_),
    .B(_14641_),
    .Y(_15641_));
 sky130_fd_sc_hd__xor2_2 _25672_ (.A(_15640_),
    .B(_15641_),
    .X(_15642_));
 sky130_fd_sc_hd__xnor2_2 _25673_ (.A(_15636_),
    .B(_15642_),
    .Y(_15644_));
 sky130_fd_sc_hd__xnor2_2 _25674_ (.A(_15635_),
    .B(_15644_),
    .Y(_15645_));
 sky130_fd_sc_hd__buf_1 _25675_ (.A(_14356_),
    .X(_15646_));
 sky130_fd_sc_hd__buf_1 _25676_ (.A(_13934_),
    .X(_15647_));
 sky130_fd_sc_hd__buf_1 _25677_ (.A(_15647_),
    .X(_15648_));
 sky130_fd_sc_hd__and4_2 _25678_ (.A(_11842_),
    .B(_12243_),
    .C(_15208_),
    .D(_14999_),
    .X(_15649_));
 sky130_fd_sc_hd__buf_1 _25679_ (.A(_13926_),
    .X(_15650_));
 sky130_fd_sc_hd__o22a_2 _25680_ (.A1(_14978_),
    .A2(_14987_),
    .B1(_15004_),
    .B2(_15650_),
    .X(_15651_));
 sky130_fd_sc_hd__o22a_2 _25681_ (.A1(_15646_),
    .A2(_15648_),
    .B1(_15649_),
    .B2(_15651_),
    .X(_15652_));
 sky130_fd_sc_hd__nor4_2 _25682_ (.A(_15646_),
    .B(_15647_),
    .C(_15649_),
    .D(_15651_),
    .Y(_15653_));
 sky130_fd_sc_hd__nor2_2 _25683_ (.A(_15652_),
    .B(_15653_),
    .Y(_15655_));
 sky130_fd_sc_hd__nor4_2 _25684_ (.A(_13844_),
    .B(_13932_),
    .C(_14364_),
    .D(_14656_),
    .Y(_15656_));
 sky130_fd_sc_hd__nor2_2 _25685_ (.A(_14993_),
    .B(_15218_),
    .Y(_15657_));
 sky130_fd_sc_hd__and3_2 _25686_ (.A(_13839_),
    .B(_15656_),
    .C(_15657_),
    .X(_15658_));
 sky130_fd_sc_hd__or2_2 _25687_ (.A(iX[11]),
    .B(iX[43]),
    .X(_15659_));
 sky130_fd_sc_hd__a32o_2 _25688_ (.A1(_15659_),
    .A2(_14365_),
    .A3(_14661_),
    .B1(_15656_),
    .B2(_13840_),
    .X(_15660_));
 sky130_fd_sc_hd__o21a_2 _25689_ (.A1(_14990_),
    .A2(_15660_),
    .B1(_15657_),
    .X(_15661_));
 sky130_fd_sc_hd__a21oi_2 _25690_ (.A1(_14991_),
    .A2(_15217_),
    .B1(_15215_),
    .Y(_15662_));
 sky130_fd_sc_hd__a211o_4 _25691_ (.A1(_13237_),
    .A2(_15658_),
    .B1(_15661_),
    .C1(_15662_),
    .X(_15663_));
 sky130_fd_sc_hd__and2_2 _25692_ (.A(iX[16]),
    .B(iX[48]),
    .X(_15664_));
 sky130_fd_sc_hd__nor2_2 _25693_ (.A(iX[16]),
    .B(iX[48]),
    .Y(_15666_));
 sky130_fd_sc_hd__nor2_2 _25694_ (.A(_15664_),
    .B(_15666_),
    .Y(_15667_));
 sky130_fd_sc_hd__xnor2_2 _25695_ (.A(_15663_),
    .B(_15667_),
    .Y(_15668_));
 sky130_fd_sc_hd__nor2_2 _25696_ (.A(_11575_),
    .B(_15668_),
    .Y(_15669_));
 sky130_fd_sc_hd__and4_2 _25697_ (.A(_11381_),
    .B(_15224_),
    .C(_15226_),
    .D(_15669_),
    .X(_15670_));
 sky130_fd_sc_hd__bufinv_8 _25698_ (.A(_15667_),
    .Y(_15671_));
 sky130_fd_sc_hd__xnor2_2 _25699_ (.A(_15663_),
    .B(_15671_),
    .Y(_15672_));
 sky130_fd_sc_hd__a32o_2 _25700_ (.A1(_11585_),
    .A2(_15224_),
    .A3(_15226_),
    .B1(_15672_),
    .B2(_11381_),
    .X(_15673_));
 sky130_fd_sc_hd__or4b_2 _25701_ (.A(_11794_),
    .B(_14998_),
    .C(_15670_),
    .D_N(_15673_),
    .X(_15674_));
 sky130_fd_sc_hd__buf_1 _25702_ (.A(_12451_),
    .X(_15675_));
 sky130_fd_sc_hd__buf_2 _25703_ (.A(_15675_),
    .X(_15677_));
 sky130_fd_sc_hd__and2_2 _25704_ (.A(_14994_),
    .B(_14996_),
    .X(_15678_));
 sky130_fd_sc_hd__buf_1 _25705_ (.A(_15678_),
    .X(_15679_));
 sky130_fd_sc_hd__or4b_2 _25706_ (.A(_11566_),
    .B(_15219_),
    .C(_15220_),
    .D_N(_15669_),
    .X(_15680_));
 sky130_fd_sc_hd__a22o_2 _25707_ (.A1(_15677_),
    .A2(_15679_),
    .B1(_15680_),
    .B2(_15673_),
    .X(_15681_));
 sky130_fd_sc_hd__a21bo_2 _25708_ (.A1(_15214_),
    .A2(_15228_),
    .B1_N(_15222_),
    .X(_15682_));
 sky130_fd_sc_hd__nand3_2 _25709_ (.A(_15674_),
    .B(_15681_),
    .C(_15682_),
    .Y(_15683_));
 sky130_fd_sc_hd__a21o_2 _25710_ (.A1(_15674_),
    .A2(_15681_),
    .B1(_15682_),
    .X(_15684_));
 sky130_fd_sc_hd__nand3_2 _25711_ (.A(_15655_),
    .B(_15683_),
    .C(_15684_),
    .Y(_15685_));
 sky130_fd_sc_hd__a21o_2 _25712_ (.A1(_15683_),
    .A2(_15684_),
    .B1(_15655_),
    .X(_15686_));
 sky130_fd_sc_hd__a21bo_2 _25713_ (.A1(_15213_),
    .A2(_15233_),
    .B1_N(_15232_),
    .X(_15688_));
 sky130_fd_sc_hd__nand3_2 _25714_ (.A(_15685_),
    .B(_15686_),
    .C(_15688_),
    .Y(_15689_));
 sky130_fd_sc_hd__a21o_2 _25715_ (.A1(_15685_),
    .A2(_15686_),
    .B1(_15688_),
    .X(_15690_));
 sky130_fd_sc_hd__nand3_2 _25716_ (.A(_15645_),
    .B(_15689_),
    .C(_15690_),
    .Y(_15691_));
 sky130_fd_sc_hd__a21o_2 _25717_ (.A1(_15689_),
    .A2(_15690_),
    .B1(_15645_),
    .X(_15692_));
 sky130_fd_sc_hd__o211ai_2 _25718_ (.A1(_15239_),
    .A2(_15241_),
    .B1(_15691_),
    .C1(_15692_),
    .Y(_15693_));
 sky130_fd_sc_hd__a211o_2 _25719_ (.A1(_15691_),
    .A2(_15692_),
    .B1(_15239_),
    .C1(_15241_),
    .X(_15694_));
 sky130_fd_sc_hd__and3_2 _25720_ (.A(_15634_),
    .B(_15693_),
    .C(_15694_),
    .X(_15695_));
 sky130_fd_sc_hd__a21oi_2 _25721_ (.A1(_15693_),
    .A2(_15694_),
    .B1(_15634_),
    .Y(_15696_));
 sky130_fd_sc_hd__a211o_2 _25722_ (.A1(_15609_),
    .A2(_15245_),
    .B1(_15695_),
    .C1(_15696_),
    .X(_15697_));
 sky130_fd_sc_hd__o211ai_2 _25723_ (.A1(_15695_),
    .A2(_15696_),
    .B1(_15609_),
    .C1(_15245_),
    .Y(_15699_));
 sky130_fd_sc_hd__nand3_2 _25724_ (.A(_15608_),
    .B(_15697_),
    .C(_15699_),
    .Y(_15700_));
 sky130_fd_sc_hd__a21o_2 _25725_ (.A1(_15697_),
    .A2(_15699_),
    .B1(_15608_),
    .X(_15701_));
 sky130_fd_sc_hd__o211ai_2 _25726_ (.A1(_15247_),
    .A2(_15582_),
    .B1(_15700_),
    .C1(_15701_),
    .Y(_15702_));
 sky130_fd_sc_hd__a211o_2 _25727_ (.A1(_15700_),
    .A2(_15701_),
    .B1(_15247_),
    .C1(_15582_),
    .X(_15703_));
 sky130_fd_sc_hd__nand3_2 _25728_ (.A(_15581_),
    .B(_15702_),
    .C(_15703_),
    .Y(_15704_));
 sky130_fd_sc_hd__a21o_2 _25729_ (.A1(_15702_),
    .A2(_15703_),
    .B1(_15581_),
    .X(_15705_));
 sky130_fd_sc_hd__nand2_2 _25730_ (.A(_15704_),
    .B(_15705_),
    .Y(_15706_));
 sky130_fd_sc_hd__xnor2_2 _25731_ (.A(_15580_),
    .B(_15706_),
    .Y(_15707_));
 sky130_fd_sc_hd__a21oi_2 _25732_ (.A1(_15262_),
    .A2(_15259_),
    .B1(_15258_),
    .Y(_15708_));
 sky130_fd_sc_hd__xnor2_2 _25733_ (.A(_15707_),
    .B(_15708_),
    .Y(_15710_));
 sky130_fd_sc_hd__xnor2_2 _25734_ (.A(_15579_),
    .B(_15710_),
    .Y(_15711_));
 sky130_fd_sc_hd__and2b_2 _25735_ (.A_N(_15122_),
    .B(_15346_),
    .X(_15712_));
 sky130_fd_sc_hd__a21o_2 _25736_ (.A1(_15266_),
    .A2(_15350_),
    .B1(_15712_),
    .X(_15713_));
 sky130_fd_sc_hd__and2b_2 _25737_ (.A_N(_15329_),
    .B(_15330_),
    .X(_15714_));
 sky130_fd_sc_hd__and2b_2 _25738_ (.A_N(_15331_),
    .B(_15338_),
    .X(_15715_));
 sky130_fd_sc_hd__or2b_2 _25739_ (.A(_15276_),
    .B_N(_15275_),
    .X(_15716_));
 sky130_fd_sc_hd__nand2_2 _25740_ (.A(_15277_),
    .B(_15283_),
    .Y(_15717_));
 sky130_fd_sc_hd__and4_2 _25741_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[45]),
    .D(iX[46]),
    .X(_15718_));
 sky130_fd_sc_hd__a22oi_2 _25742_ (.A1(iY[35]),
    .A2(iX[45]),
    .B1(iX[46]),
    .B2(iY[34]),
    .Y(_15719_));
 sky130_fd_sc_hd__nor2_2 _25743_ (.A(_15718_),
    .B(_15719_),
    .Y(_15721_));
 sky130_fd_sc_hd__nand2_2 _25744_ (.A(iY[33]),
    .B(iX[47]),
    .Y(_15722_));
 sky130_fd_sc_hd__xnor2_2 _25745_ (.A(_15721_),
    .B(_15722_),
    .Y(_15723_));
 sky130_fd_sc_hd__o21ba_2 _25746_ (.A1(_15272_),
    .A2(_15274_),
    .B1_N(_15270_),
    .X(_15724_));
 sky130_fd_sc_hd__xnor2_2 _25747_ (.A(_15723_),
    .B(_15724_),
    .Y(_15725_));
 sky130_fd_sc_hd__and4_2 _25748_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[44]),
    .D(iX[48]),
    .X(_15726_));
 sky130_fd_sc_hd__a22oi_2 _25749_ (.A1(iY[36]),
    .A2(iX[44]),
    .B1(iX[48]),
    .B2(iY[32]),
    .Y(_15727_));
 sky130_fd_sc_hd__nor2_2 _25750_ (.A(_15726_),
    .B(_15727_),
    .Y(_15728_));
 sky130_fd_sc_hd__nand2_2 _25751_ (.A(iY[37]),
    .B(iX[43]),
    .Y(_15729_));
 sky130_fd_sc_hd__xnor2_2 _25752_ (.A(_15728_),
    .B(_15729_),
    .Y(_15730_));
 sky130_fd_sc_hd__xnor2_2 _25753_ (.A(_15725_),
    .B(_15730_),
    .Y(_15732_));
 sky130_fd_sc_hd__a21o_2 _25754_ (.A1(_15716_),
    .A2(_15717_),
    .B1(_15732_),
    .X(_15733_));
 sky130_fd_sc_hd__nand3_2 _25755_ (.A(_15716_),
    .B(_15717_),
    .C(_15732_),
    .Y(_15734_));
 sky130_fd_sc_hd__o21ba_2 _25756_ (.A1(_15290_),
    .A2(_15292_),
    .B1_N(_15289_),
    .X(_15735_));
 sky130_fd_sc_hd__o21ba_2 _25757_ (.A1(_15279_),
    .A2(_15281_),
    .B1_N(_15278_),
    .X(_15736_));
 sky130_fd_sc_hd__and4_2 _25758_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[41]),
    .D(iX[42]),
    .X(_15737_));
 sky130_fd_sc_hd__a22oi_2 _25759_ (.A1(iY[39]),
    .A2(iX[41]),
    .B1(iX[42]),
    .B2(iY[38]),
    .Y(_15738_));
 sky130_fd_sc_hd__nor2_2 _25760_ (.A(_15737_),
    .B(_15738_),
    .Y(_15739_));
 sky130_fd_sc_hd__nand2_2 _25761_ (.A(iX[40]),
    .B(iY[40]),
    .Y(_15740_));
 sky130_fd_sc_hd__xnor2_2 _25762_ (.A(_15739_),
    .B(_15740_),
    .Y(_15741_));
 sky130_fd_sc_hd__xnor2_2 _25763_ (.A(_15736_),
    .B(_15741_),
    .Y(_15743_));
 sky130_fd_sc_hd__xnor2_2 _25764_ (.A(_15735_),
    .B(_15743_),
    .Y(_15744_));
 sky130_fd_sc_hd__and3_2 _25765_ (.A(_15733_),
    .B(_15734_),
    .C(_15744_),
    .X(_15745_));
 sky130_fd_sc_hd__a21oi_2 _25766_ (.A1(_15733_),
    .A2(_15734_),
    .B1(_15744_),
    .Y(_15746_));
 sky130_fd_sc_hd__or2_2 _25767_ (.A(_15745_),
    .B(_15746_),
    .X(_15747_));
 sky130_fd_sc_hd__a21o_2 _25768_ (.A1(_15285_),
    .A2(_15297_),
    .B1(_15747_),
    .X(_15748_));
 sky130_fd_sc_hd__nand3_2 _25769_ (.A(_15285_),
    .B(_15297_),
    .C(_15747_),
    .Y(_15749_));
 sky130_fd_sc_hd__and2b_2 _25770_ (.A_N(_15318_),
    .B(_15317_),
    .X(_15750_));
 sky130_fd_sc_hd__or2b_2 _25771_ (.A(_15288_),
    .B_N(_15294_),
    .X(_15751_));
 sky130_fd_sc_hd__or2b_2 _25772_ (.A(_15287_),
    .B_N(_15295_),
    .X(_15752_));
 sky130_fd_sc_hd__and4_2 _25773_ (.A(iX[35]),
    .B(iX[36]),
    .C(iY[44]),
    .D(iY[45]),
    .X(_15754_));
 sky130_fd_sc_hd__a22oi_2 _25774_ (.A1(iX[36]),
    .A2(iY[44]),
    .B1(iY[45]),
    .B2(iX[35]),
    .Y(_15755_));
 sky130_fd_sc_hd__nor2_2 _25775_ (.A(_15754_),
    .B(_15755_),
    .Y(_15756_));
 sky130_fd_sc_hd__a21oi_2 _25776_ (.A1(iX[34]),
    .A2(iY[46]),
    .B1(_15756_),
    .Y(_15757_));
 sky130_fd_sc_hd__and3_2 _25777_ (.A(iX[34]),
    .B(iY[46]),
    .C(_15756_),
    .X(_15758_));
 sky130_fd_sc_hd__nor2_2 _25778_ (.A(_15757_),
    .B(_15758_),
    .Y(_15759_));
 sky130_fd_sc_hd__and4_2 _25779_ (.A(iX[38]),
    .B(iX[39]),
    .C(iY[41]),
    .D(iY[42]),
    .X(_15760_));
 sky130_fd_sc_hd__a22oi_2 _25780_ (.A1(iX[39]),
    .A2(iY[41]),
    .B1(iY[42]),
    .B2(iX[38]),
    .Y(_15761_));
 sky130_fd_sc_hd__nor2_2 _25781_ (.A(_15760_),
    .B(_15761_),
    .Y(_15762_));
 sky130_fd_sc_hd__nand2_2 _25782_ (.A(iX[37]),
    .B(iY[43]),
    .Y(_15763_));
 sky130_fd_sc_hd__xnor2_2 _25783_ (.A(_15762_),
    .B(_15763_),
    .Y(_15765_));
 sky130_fd_sc_hd__o21ba_2 _25784_ (.A1(_15313_),
    .A2(_15316_),
    .B1_N(_15312_),
    .X(_15766_));
 sky130_fd_sc_hd__xnor2_2 _25785_ (.A(_15765_),
    .B(_15766_),
    .Y(_15767_));
 sky130_fd_sc_hd__and2_2 _25786_ (.A(_15759_),
    .B(_15767_),
    .X(_15768_));
 sky130_fd_sc_hd__nor2_2 _25787_ (.A(_15759_),
    .B(_15767_),
    .Y(_15769_));
 sky130_fd_sc_hd__or2_2 _25788_ (.A(_15768_),
    .B(_15769_),
    .X(_15770_));
 sky130_fd_sc_hd__a21o_2 _25789_ (.A1(_15751_),
    .A2(_15752_),
    .B1(_15770_),
    .X(_15771_));
 sky130_fd_sc_hd__nand3_2 _25790_ (.A(_15751_),
    .B(_15752_),
    .C(_15770_),
    .Y(_15772_));
 sky130_fd_sc_hd__o211ai_2 _25791_ (.A1(_15750_),
    .A2(_15320_),
    .B1(_15771_),
    .C1(_15772_),
    .Y(_15773_));
 sky130_fd_sc_hd__a211o_2 _25792_ (.A1(_15771_),
    .A2(_15772_),
    .B1(_15750_),
    .C1(_15320_),
    .X(_15774_));
 sky130_fd_sc_hd__nand4_2 _25793_ (.A(_15748_),
    .B(_15749_),
    .C(_15773_),
    .D(_15774_),
    .Y(_15776_));
 sky130_fd_sc_hd__a22o_2 _25794_ (.A1(_15748_),
    .A2(_15749_),
    .B1(_15773_),
    .B2(_15774_),
    .X(_15777_));
 sky130_fd_sc_hd__nand2_2 _25795_ (.A(_15776_),
    .B(_15777_),
    .Y(_15778_));
 sky130_fd_sc_hd__o21ai_2 _25796_ (.A1(_15302_),
    .A2(_15328_),
    .B1(_15300_),
    .Y(_15779_));
 sky130_fd_sc_hd__xor2_2 _25797_ (.A(_15778_),
    .B(_15779_),
    .X(_15780_));
 sky130_fd_sc_hd__nor2_2 _25798_ (.A(_15332_),
    .B(_15333_),
    .Y(_15781_));
 sky130_fd_sc_hd__a31o_2 _25799_ (.A1(iX[33]),
    .A2(iY[46]),
    .A3(_15309_),
    .B1(_15307_),
    .X(_15782_));
 sky130_fd_sc_hd__a22o_2 _25800_ (.A1(iX[33]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[32]),
    .X(_15783_));
 sky130_fd_sc_hd__nand2_2 _25801_ (.A(iX[33]),
    .B(iY[48]),
    .Y(_15784_));
 sky130_fd_sc_hd__or2_2 _25802_ (.A(_15333_),
    .B(_15784_),
    .X(_15785_));
 sky130_fd_sc_hd__nand2_2 _25803_ (.A(_15783_),
    .B(_15785_),
    .Y(_15787_));
 sky130_fd_sc_hd__xnor2_2 _25804_ (.A(_15782_),
    .B(_15787_),
    .Y(_15788_));
 sky130_fd_sc_hd__nand2_2 _25805_ (.A(_15781_),
    .B(_15788_),
    .Y(_15789_));
 sky130_fd_sc_hd__or2_2 _25806_ (.A(_15781_),
    .B(_15788_),
    .X(_15790_));
 sky130_fd_sc_hd__nand2_2 _25807_ (.A(_15789_),
    .B(_15790_),
    .Y(_15791_));
 sky130_fd_sc_hd__a21oi_2 _25808_ (.A1(_15323_),
    .A2(_15325_),
    .B1(_15791_),
    .Y(_15792_));
 sky130_fd_sc_hd__and3_2 _25809_ (.A(_15323_),
    .B(_15325_),
    .C(_15791_),
    .X(_15793_));
 sky130_fd_sc_hd__nor2_2 _25810_ (.A(_15792_),
    .B(_15793_),
    .Y(_15794_));
 sky130_fd_sc_hd__xnor2_2 _25811_ (.A(_15780_),
    .B(_15794_),
    .Y(_15795_));
 sky130_fd_sc_hd__o21ai_2 _25812_ (.A1(_15714_),
    .A2(_15715_),
    .B1(_15795_),
    .Y(_15796_));
 sky130_fd_sc_hd__or3_2 _25813_ (.A(_15714_),
    .B(_15715_),
    .C(_15795_),
    .X(_15798_));
 sky130_fd_sc_hd__nand2_2 _25814_ (.A(_15796_),
    .B(_15798_),
    .Y(_15799_));
 sky130_fd_sc_hd__xor2_2 _25815_ (.A(_15335_),
    .B(_15799_),
    .X(_15800_));
 sky130_fd_sc_hd__o21a_2 _25816_ (.A1(_15341_),
    .A2(_15343_),
    .B1(_15800_),
    .X(_15801_));
 sky130_fd_sc_hd__nor3_2 _25817_ (.A(_15341_),
    .B(_15343_),
    .C(_15800_),
    .Y(_15802_));
 sky130_fd_sc_hd__nor2_2 _25818_ (.A(_15801_),
    .B(_15802_),
    .Y(_15803_));
 sky130_fd_sc_hd__nor2_2 _25819_ (.A(_15267_),
    .B(_15345_),
    .Y(_15804_));
 sky130_fd_sc_hd__a21oi_2 _25820_ (.A1(_15347_),
    .A2(_15346_),
    .B1(_15804_),
    .Y(_15805_));
 sky130_fd_sc_hd__xnor2_2 _25821_ (.A(_15803_),
    .B(_15805_),
    .Y(_15806_));
 sky130_fd_sc_hd__xor2_2 _25822_ (.A(_15713_),
    .B(_15806_),
    .X(_15807_));
 sky130_fd_sc_hd__xor2_2 _25823_ (.A(_15711_),
    .B(_15807_),
    .X(_15809_));
 sky130_fd_sc_hd__xnor2_2 _25824_ (.A(oO[16]),
    .B(_15809_),
    .Y(_15810_));
 sky130_fd_sc_hd__and2b_2 _25825_ (.A_N(_15578_),
    .B(_15810_),
    .X(_15811_));
 sky130_fd_sc_hd__and2b_2 _25826_ (.A_N(_15810_),
    .B(_15578_),
    .X(_15812_));
 sky130_fd_sc_hd__or2_2 _25827_ (.A(_15811_),
    .B(_15812_),
    .X(_15813_));
 sky130_fd_sc_hd__a21oi_2 _25828_ (.A1(_15356_),
    .A2(_15358_),
    .B1(_15354_),
    .Y(_15814_));
 sky130_fd_sc_hd__xor2_2 _25829_ (.A(_15813_),
    .B(_15814_),
    .X(_15815_));
 sky130_fd_sc_hd__and2_2 _25830_ (.A(_15575_),
    .B(_15815_),
    .X(_15816_));
 sky130_fd_sc_hd__nor2_2 _25831_ (.A(_15575_),
    .B(_15815_),
    .Y(_15817_));
 sky130_fd_sc_hd__or2_2 _25832_ (.A(_15816_),
    .B(_15817_),
    .X(_15818_));
 sky130_fd_sc_hd__xor2_2 _25833_ (.A(_15468_),
    .B(_15818_),
    .X(oO[48]));
 sky130_fd_sc_hd__and3b_2 _25834_ (.A_N(_15258_),
    .B(_15259_),
    .C(_15262_),
    .X(_15820_));
 sky130_fd_sc_hd__a22o_2 _25835_ (.A1(_15707_),
    .A2(_15820_),
    .B1(_15710_),
    .B2(_15579_),
    .X(_15821_));
 sky130_fd_sc_hd__nand2_2 _25836_ (.A(_15258_),
    .B(_15707_),
    .Y(_15822_));
 sky130_fd_sc_hd__and3_2 _25837_ (.A(_15580_),
    .B(_15704_),
    .C(_15705_),
    .X(_15823_));
 sky130_fd_sc_hd__inv_2 _25838_ (.A(_15156_),
    .Y(_15824_));
 sky130_fd_sc_hd__nand2_2 _25839_ (.A(_15824_),
    .B(_15604_),
    .Y(_15825_));
 sky130_fd_sc_hd__and2_2 _25840_ (.A(_15612_),
    .B(_15629_),
    .X(_15826_));
 sky130_fd_sc_hd__or2_2 _25841_ (.A(_15613_),
    .B(_15614_),
    .X(_15827_));
 sky130_fd_sc_hd__or2_2 _25842_ (.A(_15615_),
    .B(_15618_),
    .X(_15828_));
 sky130_fd_sc_hd__or2_2 _25843_ (.A(iY[17]),
    .B(iY[49]),
    .X(_15830_));
 sky130_fd_sc_hd__nand2_2 _25844_ (.A(iY[17]),
    .B(iY[49]),
    .Y(_15831_));
 sky130_fd_sc_hd__nand2_2 _25845_ (.A(_15830_),
    .B(_15831_),
    .Y(_15832_));
 sky130_fd_sc_hd__a21oi_2 _25846_ (.A1(_15592_),
    .A2(_15595_),
    .B1(_15593_),
    .Y(_15833_));
 sky130_fd_sc_hd__xnor2_2 _25847_ (.A(_15832_),
    .B(_15833_),
    .Y(_15834_));
 sky130_fd_sc_hd__buf_1 _25848_ (.A(_15834_),
    .X(_15835_));
 sky130_fd_sc_hd__nor2_2 _25849_ (.A(_11578_),
    .B(_15835_),
    .Y(_15836_));
 sky130_fd_sc_hd__nor2_2 _25850_ (.A(_12468_),
    .B(_15597_),
    .Y(_15837_));
 sky130_fd_sc_hd__and3_2 _25851_ (.A(_12838_),
    .B(_15585_),
    .C(_15837_),
    .X(_15838_));
 sky130_fd_sc_hd__a21oi_2 _25852_ (.A1(_12827_),
    .A2(_15586_),
    .B1(_15600_),
    .Y(_15839_));
 sky130_fd_sc_hd__nor2_2 _25853_ (.A(_15838_),
    .B(_15839_),
    .Y(_15841_));
 sky130_fd_sc_hd__xnor2_2 _25854_ (.A(_15836_),
    .B(_15841_),
    .Y(_15842_));
 sky130_fd_sc_hd__and3_2 _25855_ (.A(_15827_),
    .B(_15828_),
    .C(_15842_),
    .X(_15843_));
 sky130_fd_sc_hd__a21oi_2 _25856_ (.A1(_15827_),
    .A2(_15828_),
    .B1(_15842_),
    .Y(_15844_));
 sky130_fd_sc_hd__nor2_2 _25857_ (.A(_15843_),
    .B(_15844_),
    .Y(_15845_));
 sky130_fd_sc_hd__o21ba_2 _25858_ (.A1(_15166_),
    .A2(_15583_),
    .B1_N(_15603_),
    .X(_15846_));
 sky130_fd_sc_hd__nor2_2 _25859_ (.A(_15601_),
    .B(_15846_),
    .Y(_15847_));
 sky130_fd_sc_hd__xnor2_2 _25860_ (.A(_15845_),
    .B(_15847_),
    .Y(_15848_));
 sky130_fd_sc_hd__o21a_2 _25861_ (.A1(_15826_),
    .A2(_15631_),
    .B1(_15848_),
    .X(_15849_));
 sky130_fd_sc_hd__or3_2 _25862_ (.A(_15826_),
    .B(_15631_),
    .C(_15848_),
    .X(_15850_));
 sky130_fd_sc_hd__and2b_2 _25863_ (.A_N(_15849_),
    .B(_15850_),
    .X(_15852_));
 sky130_fd_sc_hd__xnor2_2 _25864_ (.A(_15825_),
    .B(_15852_),
    .Y(_15853_));
 sky130_fd_sc_hd__or2_2 _25865_ (.A(_15619_),
    .B(_15628_),
    .X(_15854_));
 sky130_fd_sc_hd__o21a_2 _25866_ (.A1(_15626_),
    .A2(_15627_),
    .B1(_15854_),
    .X(_15855_));
 sky130_fd_sc_hd__and2_2 _25867_ (.A(_15636_),
    .B(_15642_),
    .X(_15856_));
 sky130_fd_sc_hd__and2b_2 _25868_ (.A_N(_15644_),
    .B(_15635_),
    .X(_15857_));
 sky130_fd_sc_hd__nand2_2 _25869_ (.A(_15624_),
    .B(_14605_),
    .Y(_15858_));
 sky130_fd_sc_hd__a22o_2 _25870_ (.A1(_12460_),
    .A2(_14410_),
    .B1(_14605_),
    .B2(_12225_),
    .X(_15859_));
 sky130_fd_sc_hd__o21a_2 _25871_ (.A1(_15614_),
    .A2(_15858_),
    .B1(_15859_),
    .X(_15860_));
 sky130_fd_sc_hd__nor2_2 _25872_ (.A(_15167_),
    .B(_14948_),
    .Y(_15861_));
 sky130_fd_sc_hd__xnor2_2 _25873_ (.A(_15860_),
    .B(_15861_),
    .Y(_15863_));
 sky130_fd_sc_hd__or4_2 _25874_ (.A(_12808_),
    .B(_13241_),
    .C(_14386_),
    .D(_13891_),
    .X(_15864_));
 sky130_fd_sc_hd__a22o_2 _25875_ (.A1(_13244_),
    .A2(_13542_),
    .B1(_13887_),
    .B2(_13501_),
    .X(_15865_));
 sky130_fd_sc_hd__nand2_2 _25876_ (.A(_15864_),
    .B(_15865_),
    .Y(_15866_));
 sky130_fd_sc_hd__nand2_2 _25877_ (.A(_12816_),
    .B(_14391_),
    .Y(_15867_));
 sky130_fd_sc_hd__xnor2_2 _25878_ (.A(_15866_),
    .B(_15867_),
    .Y(_15868_));
 sky130_fd_sc_hd__o21a_2 _25879_ (.A1(_15623_),
    .A2(_15625_),
    .B1(_15620_),
    .X(_15869_));
 sky130_fd_sc_hd__xnor2_2 _25880_ (.A(_15868_),
    .B(_15869_),
    .Y(_15870_));
 sky130_fd_sc_hd__xor2_2 _25881_ (.A(_15863_),
    .B(_15870_),
    .X(_15871_));
 sky130_fd_sc_hd__o21a_2 _25882_ (.A1(_15856_),
    .A2(_15857_),
    .B1(_15871_),
    .X(_15872_));
 sky130_fd_sc_hd__or3_2 _25883_ (.A(_15856_),
    .B(_15857_),
    .C(_15871_),
    .X(_15874_));
 sky130_fd_sc_hd__and2b_2 _25884_ (.A_N(_15872_),
    .B(_15874_),
    .X(_15875_));
 sky130_fd_sc_hd__xnor2_2 _25885_ (.A(_15855_),
    .B(_15875_),
    .Y(_15876_));
 sky130_fd_sc_hd__a21o_2 _25886_ (.A1(_15640_),
    .A2(_15641_),
    .B1(_15638_),
    .X(_15877_));
 sky130_fd_sc_hd__o22a_2 _25887_ (.A1(_12850_),
    .A2(_13842_),
    .B1(_13934_),
    .B2(_12773_),
    .X(_15878_));
 sky130_fd_sc_hd__a31o_2 _25888_ (.A1(_14637_),
    .A2(_13938_),
    .A3(_15637_),
    .B1(_15878_),
    .X(_15879_));
 sky130_fd_sc_hd__nor2_2 _25889_ (.A(_14641_),
    .B(_14983_),
    .Y(_15880_));
 sky130_fd_sc_hd__xnor2_2 _25890_ (.A(_15879_),
    .B(_15880_),
    .Y(_15881_));
 sky130_fd_sc_hd__o21a_2 _25891_ (.A1(_15649_),
    .A2(_15653_),
    .B1(_15881_),
    .X(_15882_));
 sky130_fd_sc_hd__nor3_2 _25892_ (.A(_15649_),
    .B(_15653_),
    .C(_15881_),
    .Y(_15883_));
 sky130_fd_sc_hd__or2_2 _25893_ (.A(_15882_),
    .B(_15883_),
    .X(_15885_));
 sky130_fd_sc_hd__xnor2_2 _25894_ (.A(_15877_),
    .B(_15885_),
    .Y(_15886_));
 sky130_fd_sc_hd__buf_1 _25895_ (.A(_12759_),
    .X(_15887_));
 sky130_fd_sc_hd__buf_1 _25896_ (.A(_15208_),
    .X(_15888_));
 sky130_fd_sc_hd__nand2_2 _25897_ (.A(_15887_),
    .B(_15888_),
    .Y(_15889_));
 sky130_fd_sc_hd__nand2_2 _25898_ (.A(_12243_),
    .B(_14999_),
    .Y(_15890_));
 sky130_fd_sc_hd__and3_2 _25899_ (.A(_11842_),
    .B(_14995_),
    .C(_14996_),
    .X(_15891_));
 sky130_fd_sc_hd__xnor2_2 _25900_ (.A(_15890_),
    .B(_15891_),
    .Y(_15892_));
 sky130_fd_sc_hd__xnor2_2 _25901_ (.A(_15889_),
    .B(_15892_),
    .Y(_15893_));
 sky130_fd_sc_hd__or2_2 _25902_ (.A(iX[17]),
    .B(iX[49]),
    .X(_15894_));
 sky130_fd_sc_hd__nand2_2 _25903_ (.A(iX[17]),
    .B(iX[49]),
    .Y(_15896_));
 sky130_fd_sc_hd__nand2_2 _25904_ (.A(_15894_),
    .B(_15896_),
    .Y(_15897_));
 sky130_fd_sc_hd__a21oi_2 _25905_ (.A1(_15663_),
    .A2(_15667_),
    .B1(_15664_),
    .Y(_15898_));
 sky130_fd_sc_hd__xor2_2 _25906_ (.A(_15897_),
    .B(_15898_),
    .X(_15899_));
 sky130_fd_sc_hd__buf_2 _25907_ (.A(_15899_),
    .X(_15900_));
 sky130_fd_sc_hd__and3_2 _25908_ (.A(_11380_),
    .B(_15669_),
    .C(_15900_),
    .X(_15901_));
 sky130_fd_sc_hd__a21oi_2 _25909_ (.A1(_11380_),
    .A2(_15900_),
    .B1(_15669_),
    .Y(_15902_));
 sky130_fd_sc_hd__nor2_2 _25910_ (.A(_15901_),
    .B(_15902_),
    .Y(_15903_));
 sky130_fd_sc_hd__and4_2 _25911_ (.A(_12451_),
    .B(_15223_),
    .C(_15225_),
    .D(_15903_),
    .X(_15904_));
 sky130_fd_sc_hd__a31o_2 _25912_ (.A1(_15675_),
    .A2(_15224_),
    .A3(_15226_),
    .B1(_15903_),
    .X(_15905_));
 sky130_fd_sc_hd__and2b_2 _25913_ (.A_N(_15904_),
    .B(_15905_),
    .X(_15907_));
 sky130_fd_sc_hd__a31o_2 _25914_ (.A1(_15677_),
    .A2(_15679_),
    .A3(_15673_),
    .B1(_15670_),
    .X(_15908_));
 sky130_fd_sc_hd__xor2_2 _25915_ (.A(_15907_),
    .B(_15908_),
    .X(_15909_));
 sky130_fd_sc_hd__xnor2_2 _25916_ (.A(_15893_),
    .B(_15909_),
    .Y(_15910_));
 sky130_fd_sc_hd__a21boi_2 _25917_ (.A1(_15655_),
    .A2(_15684_),
    .B1_N(_15683_),
    .Y(_15911_));
 sky130_fd_sc_hd__xor2_2 _25918_ (.A(_15910_),
    .B(_15911_),
    .X(_15912_));
 sky130_fd_sc_hd__xnor2_2 _25919_ (.A(_15886_),
    .B(_15912_),
    .Y(_15913_));
 sky130_fd_sc_hd__a21bo_2 _25920_ (.A1(_15645_),
    .A2(_15690_),
    .B1_N(_15689_),
    .X(_15914_));
 sky130_fd_sc_hd__xnor2_2 _25921_ (.A(_15913_),
    .B(_15914_),
    .Y(_15915_));
 sky130_fd_sc_hd__xor2_2 _25922_ (.A(_15876_),
    .B(_15915_),
    .X(_15916_));
 sky130_fd_sc_hd__o211a_2 _25923_ (.A1(_15239_),
    .A2(_15241_),
    .B1(_15691_),
    .C1(_15692_),
    .X(_15918_));
 sky130_fd_sc_hd__a21oi_2 _25924_ (.A1(_15634_),
    .A2(_15694_),
    .B1(_15918_),
    .Y(_15919_));
 sky130_fd_sc_hd__xnor2_2 _25925_ (.A(_15916_),
    .B(_15919_),
    .Y(_15920_));
 sky130_fd_sc_hd__xnor2_2 _25926_ (.A(_15853_),
    .B(_15920_),
    .Y(_15921_));
 sky130_fd_sc_hd__a21bo_2 _25927_ (.A1(_15608_),
    .A2(_15699_),
    .B1_N(_15697_),
    .X(_15922_));
 sky130_fd_sc_hd__xnor2_2 _25928_ (.A(_15921_),
    .B(_15922_),
    .Y(_15923_));
 sky130_fd_sc_hd__xnor2_2 _25929_ (.A(_15606_),
    .B(_15923_),
    .Y(_15924_));
 sky130_fd_sc_hd__a21boi_2 _25930_ (.A1(_15581_),
    .A2(_15703_),
    .B1_N(_15702_),
    .Y(_15925_));
 sky130_fd_sc_hd__xor2_2 _25931_ (.A(_15924_),
    .B(_15925_),
    .X(_15926_));
 sky130_fd_sc_hd__xor2_2 _25932_ (.A(_15823_),
    .B(_15926_),
    .X(_15927_));
 sky130_fd_sc_hd__xnor2_2 _25933_ (.A(_15822_),
    .B(_15927_),
    .Y(_15929_));
 sky130_fd_sc_hd__xnor2_2 _25934_ (.A(_15821_),
    .B(_15929_),
    .Y(_15930_));
 sky130_fd_sc_hd__or2b_2 _25935_ (.A(_15778_),
    .B_N(_15779_),
    .X(_15931_));
 sky130_fd_sc_hd__or3_2 _25936_ (.A(_15780_),
    .B(_15792_),
    .C(_15793_),
    .X(_15932_));
 sky130_fd_sc_hd__or2b_2 _25937_ (.A(_15724_),
    .B_N(_15723_),
    .X(_15933_));
 sky130_fd_sc_hd__nand2_2 _25938_ (.A(_15725_),
    .B(_15730_),
    .Y(_15934_));
 sky130_fd_sc_hd__and4_2 _25939_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[46]),
    .D(iX[47]),
    .X(_15935_));
 sky130_fd_sc_hd__a22oi_2 _25940_ (.A1(iY[35]),
    .A2(iX[46]),
    .B1(iX[47]),
    .B2(iY[34]),
    .Y(_15936_));
 sky130_fd_sc_hd__nor2_2 _25941_ (.A(_15935_),
    .B(_15936_),
    .Y(_15937_));
 sky130_fd_sc_hd__nand2_2 _25942_ (.A(iY[33]),
    .B(iX[48]),
    .Y(_15938_));
 sky130_fd_sc_hd__xnor2_2 _25943_ (.A(_15937_),
    .B(_15938_),
    .Y(_15940_));
 sky130_fd_sc_hd__o21ba_2 _25944_ (.A1(_15719_),
    .A2(_15722_),
    .B1_N(_15718_),
    .X(_15941_));
 sky130_fd_sc_hd__xnor2_2 _25945_ (.A(_15940_),
    .B(_15941_),
    .Y(_15942_));
 sky130_fd_sc_hd__and4_2 _25946_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[45]),
    .D(iX[49]),
    .X(_15943_));
 sky130_fd_sc_hd__a22oi_2 _25947_ (.A1(iY[36]),
    .A2(iX[45]),
    .B1(iX[49]),
    .B2(iY[32]),
    .Y(_15944_));
 sky130_fd_sc_hd__nor2_2 _25948_ (.A(_15943_),
    .B(_15944_),
    .Y(_15945_));
 sky130_fd_sc_hd__nand2_2 _25949_ (.A(iY[37]),
    .B(iX[44]),
    .Y(_15946_));
 sky130_fd_sc_hd__xnor2_2 _25950_ (.A(_15945_),
    .B(_15946_),
    .Y(_15947_));
 sky130_fd_sc_hd__xnor2_2 _25951_ (.A(_15942_),
    .B(_15947_),
    .Y(_15948_));
 sky130_fd_sc_hd__a21o_2 _25952_ (.A1(_15933_),
    .A2(_15934_),
    .B1(_15948_),
    .X(_15949_));
 sky130_fd_sc_hd__nand3_2 _25953_ (.A(_15933_),
    .B(_15934_),
    .C(_15948_),
    .Y(_15951_));
 sky130_fd_sc_hd__o21ba_2 _25954_ (.A1(_15738_),
    .A2(_15740_),
    .B1_N(_15737_),
    .X(_15952_));
 sky130_fd_sc_hd__o21ba_2 _25955_ (.A1(_15727_),
    .A2(_15729_),
    .B1_N(_15726_),
    .X(_15953_));
 sky130_fd_sc_hd__and4_2 _25956_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[42]),
    .D(iX[43]),
    .X(_15954_));
 sky130_fd_sc_hd__a22oi_2 _25957_ (.A1(iY[39]),
    .A2(iX[42]),
    .B1(iX[43]),
    .B2(iY[38]),
    .Y(_15955_));
 sky130_fd_sc_hd__nor2_2 _25958_ (.A(_15954_),
    .B(_15955_),
    .Y(_15956_));
 sky130_fd_sc_hd__nand2_2 _25959_ (.A(iY[40]),
    .B(iX[41]),
    .Y(_15957_));
 sky130_fd_sc_hd__xnor2_2 _25960_ (.A(_15956_),
    .B(_15957_),
    .Y(_15958_));
 sky130_fd_sc_hd__xnor2_2 _25961_ (.A(_15953_),
    .B(_15958_),
    .Y(_15959_));
 sky130_fd_sc_hd__xnor2_2 _25962_ (.A(_15952_),
    .B(_15959_),
    .Y(_15960_));
 sky130_fd_sc_hd__nand3_2 _25963_ (.A(_15949_),
    .B(_15951_),
    .C(_15960_),
    .Y(_15962_));
 sky130_fd_sc_hd__a21o_2 _25964_ (.A1(_15949_),
    .A2(_15951_),
    .B1(_15960_),
    .X(_15963_));
 sky130_fd_sc_hd__a21bo_2 _25965_ (.A1(_15734_),
    .A2(_15744_),
    .B1_N(_15733_),
    .X(_15964_));
 sky130_fd_sc_hd__and3_2 _25966_ (.A(_15962_),
    .B(_15963_),
    .C(_15964_),
    .X(_15965_));
 sky130_fd_sc_hd__a21oi_2 _25967_ (.A1(_15962_),
    .A2(_15963_),
    .B1(_15964_),
    .Y(_15966_));
 sky130_fd_sc_hd__nor2_2 _25968_ (.A(_15965_),
    .B(_15966_),
    .Y(_15967_));
 sky130_fd_sc_hd__and2b_2 _25969_ (.A_N(_15766_),
    .B(_15765_),
    .X(_15968_));
 sky130_fd_sc_hd__or2b_2 _25970_ (.A(_15736_),
    .B_N(_15741_),
    .X(_15969_));
 sky130_fd_sc_hd__or2b_2 _25971_ (.A(_15735_),
    .B_N(_15743_),
    .X(_15970_));
 sky130_fd_sc_hd__and4_2 _25972_ (.A(iX[36]),
    .B(iX[37]),
    .C(iY[44]),
    .D(iY[45]),
    .X(_15971_));
 sky130_fd_sc_hd__a22oi_2 _25973_ (.A1(iX[37]),
    .A2(iY[44]),
    .B1(iY[45]),
    .B2(iX[36]),
    .Y(_15973_));
 sky130_fd_sc_hd__nor2_2 _25974_ (.A(_15971_),
    .B(_15973_),
    .Y(_15974_));
 sky130_fd_sc_hd__nand2_2 _25975_ (.A(iX[35]),
    .B(iY[46]),
    .Y(_15975_));
 sky130_fd_sc_hd__xnor2_2 _25976_ (.A(_15974_),
    .B(_15975_),
    .Y(_15976_));
 sky130_fd_sc_hd__and4_2 _25977_ (.A(iX[39]),
    .B(iX[40]),
    .C(iY[41]),
    .D(iY[42]),
    .X(_15977_));
 sky130_fd_sc_hd__a22oi_2 _25978_ (.A1(iX[40]),
    .A2(iY[41]),
    .B1(iY[42]),
    .B2(iX[39]),
    .Y(_15978_));
 sky130_fd_sc_hd__nor2_2 _25979_ (.A(_15977_),
    .B(_15978_),
    .Y(_15979_));
 sky130_fd_sc_hd__nand2_2 _25980_ (.A(iX[38]),
    .B(iY[43]),
    .Y(_15980_));
 sky130_fd_sc_hd__xnor2_2 _25981_ (.A(_15979_),
    .B(_15980_),
    .Y(_15981_));
 sky130_fd_sc_hd__o21ba_2 _25982_ (.A1(_15761_),
    .A2(_15763_),
    .B1_N(_15760_),
    .X(_15982_));
 sky130_fd_sc_hd__xnor2_2 _25983_ (.A(_15981_),
    .B(_15982_),
    .Y(_15984_));
 sky130_fd_sc_hd__and2_2 _25984_ (.A(_15976_),
    .B(_15984_),
    .X(_15985_));
 sky130_fd_sc_hd__nor2_2 _25985_ (.A(_15976_),
    .B(_15984_),
    .Y(_15986_));
 sky130_fd_sc_hd__or2_2 _25986_ (.A(_15985_),
    .B(_15986_),
    .X(_15987_));
 sky130_fd_sc_hd__a21o_2 _25987_ (.A1(_15969_),
    .A2(_15970_),
    .B1(_15987_),
    .X(_15988_));
 sky130_fd_sc_hd__nand3_2 _25988_ (.A(_15969_),
    .B(_15970_),
    .C(_15987_),
    .Y(_15989_));
 sky130_fd_sc_hd__o211ai_2 _25989_ (.A1(_15968_),
    .A2(_15768_),
    .B1(_15988_),
    .C1(_15989_),
    .Y(_15990_));
 sky130_fd_sc_hd__a211o_2 _25990_ (.A1(_15988_),
    .A2(_15989_),
    .B1(_15968_),
    .C1(_15768_),
    .X(_15991_));
 sky130_fd_sc_hd__and3_2 _25991_ (.A(_15967_),
    .B(_15990_),
    .C(_15991_),
    .X(_15992_));
 sky130_fd_sc_hd__a21oi_2 _25992_ (.A1(_15990_),
    .A2(_15991_),
    .B1(_15967_),
    .Y(_15993_));
 sky130_fd_sc_hd__a211o_2 _25993_ (.A1(_15748_),
    .A2(_15776_),
    .B1(_15992_),
    .C1(_15993_),
    .X(_15995_));
 sky130_fd_sc_hd__o211ai_2 _25994_ (.A1(_15992_),
    .A2(_15993_),
    .B1(_15748_),
    .C1(_15776_),
    .Y(_15996_));
 sky130_fd_sc_hd__nand2_2 _25995_ (.A(iX[34]),
    .B(iY[47]),
    .Y(_15997_));
 sky130_fd_sc_hd__and4_2 _25996_ (.A(iX[33]),
    .B(iX[34]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_15998_));
 sky130_fd_sc_hd__a21oi_2 _25997_ (.A1(_15784_),
    .A2(_15997_),
    .B1(_15998_),
    .Y(_15999_));
 sky130_fd_sc_hd__nand2_2 _25998_ (.A(iX[32]),
    .B(iY[49]),
    .Y(_16000_));
 sky130_fd_sc_hd__xnor2_2 _25999_ (.A(_15999_),
    .B(_16000_),
    .Y(_16001_));
 sky130_fd_sc_hd__nor3_2 _26000_ (.A(_15754_),
    .B(_15758_),
    .C(_16001_),
    .Y(_16002_));
 sky130_fd_sc_hd__o21a_2 _26001_ (.A1(_15754_),
    .A2(_15758_),
    .B1(_16001_),
    .X(_16003_));
 sky130_fd_sc_hd__nor2_2 _26002_ (.A(_16002_),
    .B(_16003_),
    .Y(_16004_));
 sky130_fd_sc_hd__nor2_2 _26003_ (.A(_15333_),
    .B(_15784_),
    .Y(_16006_));
 sky130_fd_sc_hd__and3_2 _26004_ (.A(_15782_),
    .B(_15783_),
    .C(_15785_),
    .X(_16007_));
 sky130_fd_sc_hd__or2_2 _26005_ (.A(_16006_),
    .B(_16007_),
    .X(_16008_));
 sky130_fd_sc_hd__xnor2_2 _26006_ (.A(_16004_),
    .B(_16008_),
    .Y(_16009_));
 sky130_fd_sc_hd__a21o_2 _26007_ (.A1(_15771_),
    .A2(_15773_),
    .B1(_16009_),
    .X(_16010_));
 sky130_fd_sc_hd__nand3_2 _26008_ (.A(_15771_),
    .B(_15773_),
    .C(_16009_),
    .Y(_16011_));
 sky130_fd_sc_hd__nand2_2 _26009_ (.A(_16010_),
    .B(_16011_),
    .Y(_16012_));
 sky130_fd_sc_hd__xor2_2 _26010_ (.A(_15789_),
    .B(_16012_),
    .X(_16013_));
 sky130_fd_sc_hd__a21oi_2 _26011_ (.A1(_15995_),
    .A2(_15996_),
    .B1(_16013_),
    .Y(_16014_));
 sky130_fd_sc_hd__and3_2 _26012_ (.A(_15995_),
    .B(_15996_),
    .C(_16013_),
    .X(_16015_));
 sky130_fd_sc_hd__a211o_2 _26013_ (.A1(_15931_),
    .A2(_15932_),
    .B1(_16014_),
    .C1(_16015_),
    .X(_16017_));
 sky130_fd_sc_hd__o211ai_2 _26014_ (.A1(_16014_),
    .A2(_16015_),
    .B1(_15931_),
    .C1(_15932_),
    .Y(_16018_));
 sky130_fd_sc_hd__and3_2 _26015_ (.A(_15792_),
    .B(_16017_),
    .C(_16018_),
    .X(_16019_));
 sky130_fd_sc_hd__a21oi_2 _26016_ (.A1(_16017_),
    .A2(_16018_),
    .B1(_15792_),
    .Y(_16020_));
 sky130_fd_sc_hd__nor2_2 _26017_ (.A(_16019_),
    .B(_16020_),
    .Y(_16021_));
 sky130_fd_sc_hd__o21a_2 _26018_ (.A1(_15335_),
    .A2(_15799_),
    .B1(_15796_),
    .X(_16022_));
 sky130_fd_sc_hd__xnor2_2 _26019_ (.A(_16021_),
    .B(_16022_),
    .Y(_16023_));
 sky130_fd_sc_hd__and2_2 _26020_ (.A(_15801_),
    .B(_16023_),
    .X(_16024_));
 sky130_fd_sc_hd__nor2_2 _26021_ (.A(_15801_),
    .B(_16023_),
    .Y(_16025_));
 sky130_fd_sc_hd__nor2_2 _26022_ (.A(_16024_),
    .B(_16025_),
    .Y(_16026_));
 sky130_fd_sc_hd__a21o_2 _26023_ (.A1(_15804_),
    .A2(_15803_),
    .B1(_16026_),
    .X(_16028_));
 sky130_fd_sc_hd__and3_2 _26024_ (.A(_15804_),
    .B(_15803_),
    .C(_16026_),
    .X(_16029_));
 sky130_fd_sc_hd__inv_2 _26025_ (.A(_16029_),
    .Y(_16030_));
 sky130_fd_sc_hd__nand2_2 _26026_ (.A(_16028_),
    .B(_16030_),
    .Y(_16031_));
 sky130_fd_sc_hd__and3_2 _26027_ (.A(_15347_),
    .B(_15346_),
    .C(_15803_),
    .X(_16032_));
 sky130_fd_sc_hd__a21oi_2 _26028_ (.A1(_15713_),
    .A2(_15806_),
    .B1(_16032_),
    .Y(_16033_));
 sky130_fd_sc_hd__xnor2_2 _26029_ (.A(_16031_),
    .B(_16033_),
    .Y(_16034_));
 sky130_fd_sc_hd__xnor2_2 _26030_ (.A(_15930_),
    .B(_16034_),
    .Y(_16035_));
 sky130_fd_sc_hd__xor2_2 _26031_ (.A(oO[17]),
    .B(_16035_),
    .X(_16036_));
 sky130_fd_sc_hd__or2_2 _26032_ (.A(_15711_),
    .B(_15807_),
    .X(_16037_));
 sky130_fd_sc_hd__or2b_2 _26033_ (.A(oO[16]),
    .B_N(_15809_),
    .X(_16039_));
 sky130_fd_sc_hd__nand2_2 _26034_ (.A(_16037_),
    .B(_16039_),
    .Y(_16040_));
 sky130_fd_sc_hd__xor2_2 _26035_ (.A(_16036_),
    .B(_16040_),
    .X(_16041_));
 sky130_fd_sc_hd__o21ba_2 _26036_ (.A1(_15813_),
    .A2(_15814_),
    .B1_N(_15811_),
    .X(_16042_));
 sky130_fd_sc_hd__xnor2_2 _26037_ (.A(_16041_),
    .B(_16042_),
    .Y(_16043_));
 sky130_fd_sc_hd__and4_2 _26038_ (.A(iY[21]),
    .B(iY[22]),
    .C(iX[27]),
    .D(iX[28]),
    .X(_16044_));
 sky130_fd_sc_hd__a22oi_2 _26039_ (.A1(iY[22]),
    .A2(iX[27]),
    .B1(iX[28]),
    .B2(iY[21]),
    .Y(_16045_));
 sky130_fd_sc_hd__or2_2 _26040_ (.A(_16044_),
    .B(_16045_),
    .X(_16046_));
 sky130_fd_sc_hd__nand2_2 _26041_ (.A(iY[23]),
    .B(iX[26]),
    .Y(_16047_));
 sky130_fd_sc_hd__nor2_2 _26042_ (.A(_16046_),
    .B(_16047_),
    .Y(_16048_));
 sky130_fd_sc_hd__and2_2 _26043_ (.A(_16046_),
    .B(_16047_),
    .X(_16050_));
 sky130_fd_sc_hd__nor2_2 _26044_ (.A(_16048_),
    .B(_16050_),
    .Y(_16051_));
 sky130_fd_sc_hd__inv_2 _26045_ (.A(_16051_),
    .Y(_16052_));
 sky130_fd_sc_hd__a21o_2 _26046_ (.A1(iY[18]),
    .A2(iX[31]),
    .B1(_15487_),
    .X(_16053_));
 sky130_fd_sc_hd__inv_2 _26047_ (.A(_16053_),
    .Y(_16054_));
 sky130_fd_sc_hd__and3_2 _26048_ (.A(iY[18]),
    .B(iX[31]),
    .C(_15487_),
    .X(_16055_));
 sky130_fd_sc_hd__nor2_2 _26049_ (.A(_16054_),
    .B(_16055_),
    .Y(_16056_));
 sky130_fd_sc_hd__nand2_2 _26050_ (.A(iY[20]),
    .B(iX[29]),
    .Y(_16057_));
 sky130_fd_sc_hd__xnor2_2 _26051_ (.A(_16056_),
    .B(_16057_),
    .Y(_16058_));
 sky130_fd_sc_hd__o21ba_2 _26052_ (.A1(_15490_),
    .A2(_15492_),
    .B1_N(_15488_),
    .X(_16059_));
 sky130_fd_sc_hd__xor2_2 _26053_ (.A(_16058_),
    .B(_16059_),
    .X(_16061_));
 sky130_fd_sc_hd__nor2_2 _26054_ (.A(_16052_),
    .B(_16061_),
    .Y(_16062_));
 sky130_fd_sc_hd__and2_2 _26055_ (.A(_16052_),
    .B(_16061_),
    .X(_16063_));
 sky130_fd_sc_hd__or2_2 _26056_ (.A(_16062_),
    .B(_16063_),
    .X(_16064_));
 sky130_fd_sc_hd__or3_2 _26057_ (.A(_15364_),
    .B(_15365_),
    .C(_16064_),
    .X(_16065_));
 sky130_fd_sc_hd__o21ai_2 _26058_ (.A1(_15364_),
    .A2(_15365_),
    .B1(_16064_),
    .Y(_16066_));
 sky130_fd_sc_hd__nand2_2 _26059_ (.A(_16065_),
    .B(_16066_),
    .Y(_16067_));
 sky130_fd_sc_hd__a31o_2 _26060_ (.A1(_15367_),
    .A2(_15368_),
    .A3(_15480_),
    .B1(_15499_),
    .X(_16068_));
 sky130_fd_sc_hd__and2b_2 _26061_ (.A_N(_16067_),
    .B(_16068_),
    .X(_16069_));
 sky130_fd_sc_hd__and2b_2 _26062_ (.A_N(_16068_),
    .B(_16067_),
    .X(_16070_));
 sky130_fd_sc_hd__or2_2 _26063_ (.A(_16069_),
    .B(_16070_),
    .X(_16072_));
 sky130_fd_sc_hd__inv_2 _26064_ (.A(_15543_),
    .Y(_16073_));
 sky130_fd_sc_hd__or2b_2 _26065_ (.A(_15512_),
    .B_N(_15510_),
    .X(_16074_));
 sky130_fd_sc_hd__and4_2 _26066_ (.A(iX[21]),
    .B(iX[22]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_16075_));
 sky130_fd_sc_hd__a22oi_2 _26067_ (.A1(iX[22]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[21]),
    .Y(_16076_));
 sky130_fd_sc_hd__nor2_2 _26068_ (.A(_16075_),
    .B(_16076_),
    .Y(_16077_));
 sky130_fd_sc_hd__nand2_2 _26069_ (.A(iX[20]),
    .B(iY[29]),
    .Y(_16078_));
 sky130_fd_sc_hd__xnor2_2 _26070_ (.A(_16077_),
    .B(_16078_),
    .Y(_16079_));
 sky130_fd_sc_hd__o21ba_2 _26071_ (.A1(_15507_),
    .A2(_15509_),
    .B1_N(_15506_),
    .X(_16080_));
 sky130_fd_sc_hd__xnor2_2 _26072_ (.A(_16079_),
    .B(_16080_),
    .Y(_16081_));
 sky130_fd_sc_hd__nand3_2 _26073_ (.A(iX[19]),
    .B(iY[30]),
    .C(_16081_),
    .Y(_16083_));
 sky130_fd_sc_hd__a21o_2 _26074_ (.A1(iX[19]),
    .A2(iY[30]),
    .B1(_16081_),
    .X(_16084_));
 sky130_fd_sc_hd__nand2_2 _26075_ (.A(_16083_),
    .B(_16084_),
    .Y(_16085_));
 sky130_fd_sc_hd__a21oi_2 _26076_ (.A1(_16074_),
    .A2(_15514_),
    .B1(_16085_),
    .Y(_16086_));
 sky130_fd_sc_hd__and3_2 _26077_ (.A(_16074_),
    .B(_15514_),
    .C(_16085_),
    .X(_16087_));
 sky130_fd_sc_hd__nor2_2 _26078_ (.A(_16086_),
    .B(_16087_),
    .Y(_16088_));
 sky130_fd_sc_hd__nand2_2 _26079_ (.A(iX[18]),
    .B(iY[31]),
    .Y(_16089_));
 sky130_fd_sc_hd__xnor2_2 _26080_ (.A(_16088_),
    .B(_16089_),
    .Y(_16090_));
 sky130_fd_sc_hd__or2b_2 _26081_ (.A(_15529_),
    .B_N(_15535_),
    .X(_16091_));
 sky130_fd_sc_hd__or2b_2 _26082_ (.A(_15528_),
    .B_N(_15536_),
    .X(_16092_));
 sky130_fd_sc_hd__and2b_2 _26083_ (.A_N(_15494_),
    .B(_15493_),
    .X(_16093_));
 sky130_fd_sc_hd__o21ba_2 _26084_ (.A1(_15531_),
    .A2(_15534_),
    .B1_N(_15530_),
    .X(_16094_));
 sky130_fd_sc_hd__o21ba_2 _26085_ (.A1(_15483_),
    .A2(_15485_),
    .B1_N(_15482_),
    .X(_16095_));
 sky130_fd_sc_hd__and4_2 _26086_ (.A(iX[24]),
    .B(iY[24]),
    .C(iX[25]),
    .D(iY[25]),
    .X(_16096_));
 sky130_fd_sc_hd__a22oi_2 _26087_ (.A1(iY[24]),
    .A2(iX[25]),
    .B1(iY[25]),
    .B2(iX[24]),
    .Y(_16097_));
 sky130_fd_sc_hd__nor2_2 _26088_ (.A(_16096_),
    .B(_16097_),
    .Y(_16098_));
 sky130_fd_sc_hd__nand2_2 _26089_ (.A(iX[23]),
    .B(iY[26]),
    .Y(_16099_));
 sky130_fd_sc_hd__xnor2_2 _26090_ (.A(_16098_),
    .B(_16099_),
    .Y(_16100_));
 sky130_fd_sc_hd__xnor2_2 _26091_ (.A(_16095_),
    .B(_16100_),
    .Y(_16101_));
 sky130_fd_sc_hd__xnor2_2 _26092_ (.A(_16094_),
    .B(_16101_),
    .Y(_16102_));
 sky130_fd_sc_hd__o21a_2 _26093_ (.A1(_16093_),
    .A2(_15496_),
    .B1(_16102_),
    .X(_16104_));
 sky130_fd_sc_hd__nor3_2 _26094_ (.A(_16093_),
    .B(_15496_),
    .C(_16102_),
    .Y(_16105_));
 sky130_fd_sc_hd__a211oi_2 _26095_ (.A1(_16091_),
    .A2(_16092_),
    .B1(_16104_),
    .C1(_16105_),
    .Y(_16106_));
 sky130_fd_sc_hd__o211a_2 _26096_ (.A1(_16104_),
    .A2(_16105_),
    .B1(_16091_),
    .C1(_16092_),
    .X(_16107_));
 sky130_fd_sc_hd__nor2_2 _26097_ (.A(_15538_),
    .B(_15540_),
    .Y(_16108_));
 sky130_fd_sc_hd__or3_2 _26098_ (.A(_16106_),
    .B(_16107_),
    .C(_16108_),
    .X(_16109_));
 sky130_fd_sc_hd__o21ai_2 _26099_ (.A1(_16106_),
    .A2(_16107_),
    .B1(_16108_),
    .Y(_16110_));
 sky130_fd_sc_hd__and3_2 _26100_ (.A(_16090_),
    .B(_16109_),
    .C(_16110_),
    .X(_16111_));
 sky130_fd_sc_hd__a21oi_2 _26101_ (.A1(_16109_),
    .A2(_16110_),
    .B1(_16090_),
    .Y(_16112_));
 sky130_fd_sc_hd__or3_2 _26102_ (.A(_15502_),
    .B(_16111_),
    .C(_16112_),
    .X(_16113_));
 sky130_fd_sc_hd__o21ai_2 _26103_ (.A1(_16111_),
    .A2(_16112_),
    .B1(_15502_),
    .Y(_16115_));
 sky130_fd_sc_hd__o211a_2 _26104_ (.A1(_16073_),
    .A2(_15546_),
    .B1(_16113_),
    .C1(_16115_),
    .X(_16116_));
 sky130_fd_sc_hd__a211oi_2 _26105_ (.A1(_16113_),
    .A2(_16115_),
    .B1(_16073_),
    .C1(_15546_),
    .Y(_16117_));
 sky130_fd_sc_hd__or3_2 _26106_ (.A(_16072_),
    .B(_16116_),
    .C(_16117_),
    .X(_16118_));
 sky130_fd_sc_hd__o21ai_2 _26107_ (.A1(_16116_),
    .A2(_16117_),
    .B1(_16072_),
    .Y(_16119_));
 sky130_fd_sc_hd__and3_2 _26108_ (.A(_15553_),
    .B(_16118_),
    .C(_16119_),
    .X(_16120_));
 sky130_fd_sc_hd__a21oi_2 _26109_ (.A1(_16118_),
    .A2(_16119_),
    .B1(_15553_),
    .Y(_16121_));
 sky130_fd_sc_hd__a211oi_2 _26110_ (.A1(_15548_),
    .A2(_15551_),
    .B1(_16120_),
    .C1(_16121_),
    .Y(_16122_));
 sky130_fd_sc_hd__o211a_2 _26111_ (.A1(_16120_),
    .A2(_16121_),
    .B1(_15548_),
    .C1(_15551_),
    .X(_16123_));
 sky130_fd_sc_hd__a211oi_2 _26112_ (.A1(_15556_),
    .A2(_15558_),
    .B1(_16122_),
    .C1(_16123_),
    .Y(_16124_));
 sky130_fd_sc_hd__o211a_2 _26113_ (.A1(_16122_),
    .A2(_16123_),
    .B1(_15556_),
    .C1(_15558_),
    .X(_16126_));
 sky130_fd_sc_hd__a211oi_2 _26114_ (.A1(_15517_),
    .A2(_15523_),
    .B1(_16124_),
    .C1(_16126_),
    .Y(_16127_));
 sky130_fd_sc_hd__o211a_2 _26115_ (.A1(_16124_),
    .A2(_16126_),
    .B1(_15517_),
    .C1(_15523_),
    .X(_16128_));
 sky130_fd_sc_hd__o211ai_2 _26116_ (.A1(_16127_),
    .A2(_16128_),
    .B1(_15562_),
    .C1(_15565_),
    .Y(_16129_));
 sky130_fd_sc_hd__inv_2 _26117_ (.A(_16129_),
    .Y(_16130_));
 sky130_fd_sc_hd__a211oi_2 _26118_ (.A1(_15562_),
    .A2(_15565_),
    .B1(_16127_),
    .C1(_16128_),
    .Y(_16131_));
 sky130_fd_sc_hd__nor2_2 _26119_ (.A(_16130_),
    .B(_16131_),
    .Y(_16132_));
 sky130_fd_sc_hd__a21oi_2 _26120_ (.A1(_15477_),
    .A2(_15572_),
    .B1(_15570_),
    .Y(_16133_));
 sky130_fd_sc_hd__xor2_2 _26121_ (.A(_16132_),
    .B(_16133_),
    .X(_16134_));
 sky130_fd_sc_hd__nor2_2 _26122_ (.A(_16043_),
    .B(_16134_),
    .Y(_16135_));
 sky130_fd_sc_hd__nand2_2 _26123_ (.A(_16043_),
    .B(_16134_),
    .Y(_16137_));
 sky130_fd_sc_hd__or2b_2 _26124_ (.A(_16135_),
    .B_N(_16137_),
    .X(_16138_));
 sky130_fd_sc_hd__o21bai_2 _26125_ (.A1(_15468_),
    .A2(_15818_),
    .B1_N(_15816_),
    .Y(_16139_));
 sky130_fd_sc_hd__xnor2_2 _26126_ (.A(_16138_),
    .B(_16139_),
    .Y(oO[49]));
 sky130_fd_sc_hd__o21ba_2 _26127_ (.A1(_16087_),
    .A2(_16089_),
    .B1_N(_16086_),
    .X(_16140_));
 sky130_fd_sc_hd__inv_2 _26128_ (.A(_16113_),
    .Y(_16141_));
 sky130_fd_sc_hd__and3_2 _26129_ (.A(iY[20]),
    .B(iX[31]),
    .C(_15487_),
    .X(_16142_));
 sky130_fd_sc_hd__a22oi_2 _26130_ (.A1(iY[20]),
    .A2(iX[30]),
    .B1(iX[31]),
    .B2(iY[19]),
    .Y(_16143_));
 sky130_fd_sc_hd__or2_2 _26131_ (.A(_16142_),
    .B(_16143_),
    .X(_16144_));
 sky130_fd_sc_hd__a31o_2 _26132_ (.A1(iY[20]),
    .A2(iX[29]),
    .A3(_16053_),
    .B1(_16055_),
    .X(_16145_));
 sky130_fd_sc_hd__xnor2_2 _26133_ (.A(_16144_),
    .B(_16145_),
    .Y(_16147_));
 sky130_fd_sc_hd__and4_2 _26134_ (.A(iY[21]),
    .B(iY[22]),
    .C(iX[28]),
    .D(iX[29]),
    .X(_16148_));
 sky130_fd_sc_hd__a22oi_2 _26135_ (.A1(iY[22]),
    .A2(iX[28]),
    .B1(iX[29]),
    .B2(iY[21]),
    .Y(_16149_));
 sky130_fd_sc_hd__nor2_2 _26136_ (.A(_16148_),
    .B(_16149_),
    .Y(_16150_));
 sky130_fd_sc_hd__nand2_2 _26137_ (.A(iY[23]),
    .B(iX[27]),
    .Y(_16151_));
 sky130_fd_sc_hd__xnor2_2 _26138_ (.A(_16150_),
    .B(_16151_),
    .Y(_16152_));
 sky130_fd_sc_hd__nand2_2 _26139_ (.A(_16147_),
    .B(_16152_),
    .Y(_16153_));
 sky130_fd_sc_hd__or2_2 _26140_ (.A(_16147_),
    .B(_16152_),
    .X(_16154_));
 sky130_fd_sc_hd__nand2_2 _26141_ (.A(_16153_),
    .B(_16154_),
    .Y(_16155_));
 sky130_fd_sc_hd__or2_2 _26142_ (.A(_16065_),
    .B(_16155_),
    .X(_16156_));
 sky130_fd_sc_hd__nand2_2 _26143_ (.A(_16065_),
    .B(_16155_),
    .Y(_16158_));
 sky130_fd_sc_hd__nand2_2 _26144_ (.A(_16156_),
    .B(_16158_),
    .Y(_16159_));
 sky130_fd_sc_hd__inv_2 _26145_ (.A(_16111_),
    .Y(_16160_));
 sky130_fd_sc_hd__or2b_2 _26146_ (.A(_16080_),
    .B_N(_16079_),
    .X(_16161_));
 sky130_fd_sc_hd__and4_2 _26147_ (.A(iX[22]),
    .B(iX[23]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_16162_));
 sky130_fd_sc_hd__a22oi_2 _26148_ (.A1(iX[23]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[22]),
    .Y(_16163_));
 sky130_fd_sc_hd__nor2_2 _26149_ (.A(_16162_),
    .B(_16163_),
    .Y(_16164_));
 sky130_fd_sc_hd__nand2_2 _26150_ (.A(iX[21]),
    .B(iY[29]),
    .Y(_16165_));
 sky130_fd_sc_hd__xnor2_2 _26151_ (.A(_16164_),
    .B(_16165_),
    .Y(_16166_));
 sky130_fd_sc_hd__o21ba_2 _26152_ (.A1(_16076_),
    .A2(_16078_),
    .B1_N(_16075_),
    .X(_16167_));
 sky130_fd_sc_hd__xnor2_2 _26153_ (.A(_16166_),
    .B(_16167_),
    .Y(_16169_));
 sky130_fd_sc_hd__and2_2 _26154_ (.A(iX[20]),
    .B(iY[30]),
    .X(_16170_));
 sky130_fd_sc_hd__or2_2 _26155_ (.A(_16169_),
    .B(_16170_),
    .X(_16171_));
 sky130_fd_sc_hd__nand2_2 _26156_ (.A(_16169_),
    .B(_16170_),
    .Y(_16172_));
 sky130_fd_sc_hd__nand2_2 _26157_ (.A(_16171_),
    .B(_16172_),
    .Y(_16173_));
 sky130_fd_sc_hd__a21oi_2 _26158_ (.A1(_16161_),
    .A2(_16083_),
    .B1(_16173_),
    .Y(_16174_));
 sky130_fd_sc_hd__and3_2 _26159_ (.A(_16161_),
    .B(_16083_),
    .C(_16173_),
    .X(_16175_));
 sky130_fd_sc_hd__nor2_2 _26160_ (.A(_16174_),
    .B(_16175_),
    .Y(_16176_));
 sky130_fd_sc_hd__nand2_2 _26161_ (.A(iX[19]),
    .B(iY[31]),
    .Y(_16177_));
 sky130_fd_sc_hd__xnor2_2 _26162_ (.A(_16176_),
    .B(_16177_),
    .Y(_16178_));
 sky130_fd_sc_hd__or2b_2 _26163_ (.A(_16095_),
    .B_N(_16100_),
    .X(_16180_));
 sky130_fd_sc_hd__or2b_2 _26164_ (.A(_16094_),
    .B_N(_16101_),
    .X(_16181_));
 sky130_fd_sc_hd__and2b_2 _26165_ (.A_N(_16059_),
    .B(_16058_),
    .X(_16182_));
 sky130_fd_sc_hd__o21ba_2 _26166_ (.A1(_16097_),
    .A2(_16099_),
    .B1_N(_16096_),
    .X(_16183_));
 sky130_fd_sc_hd__and4_2 _26167_ (.A(iY[24]),
    .B(iX[25]),
    .C(iY[25]),
    .D(iX[26]),
    .X(_16184_));
 sky130_fd_sc_hd__a22oi_2 _26168_ (.A1(iX[25]),
    .A2(iY[25]),
    .B1(iX[26]),
    .B2(iY[24]),
    .Y(_16185_));
 sky130_fd_sc_hd__and4bb_2 _26169_ (.A_N(_16184_),
    .B_N(_16185_),
    .C(iX[24]),
    .D(iY[26]),
    .X(_16186_));
 sky130_fd_sc_hd__o2bb2a_2 _26170_ (.A1_N(iX[24]),
    .A2_N(iY[26]),
    .B1(_16184_),
    .B2(_16185_),
    .X(_16187_));
 sky130_fd_sc_hd__nor2_2 _26171_ (.A(_16186_),
    .B(_16187_),
    .Y(_16188_));
 sky130_fd_sc_hd__o21ai_2 _26172_ (.A1(_16044_),
    .A2(_16048_),
    .B1(_16188_),
    .Y(_16189_));
 sky130_fd_sc_hd__or3_2 _26173_ (.A(_16044_),
    .B(_16048_),
    .C(_16188_),
    .X(_16191_));
 sky130_fd_sc_hd__and2_2 _26174_ (.A(_16189_),
    .B(_16191_),
    .X(_16192_));
 sky130_fd_sc_hd__xnor2_2 _26175_ (.A(_16183_),
    .B(_16192_),
    .Y(_16193_));
 sky130_fd_sc_hd__o21a_2 _26176_ (.A1(_16182_),
    .A2(_16062_),
    .B1(_16193_),
    .X(_16194_));
 sky130_fd_sc_hd__nor3_2 _26177_ (.A(_16182_),
    .B(_16062_),
    .C(_16193_),
    .Y(_16195_));
 sky130_fd_sc_hd__a211oi_2 _26178_ (.A1(_16180_),
    .A2(_16181_),
    .B1(_16194_),
    .C1(_16195_),
    .Y(_16196_));
 sky130_fd_sc_hd__o211a_2 _26179_ (.A1(_16194_),
    .A2(_16195_),
    .B1(_16180_),
    .C1(_16181_),
    .X(_16197_));
 sky130_fd_sc_hd__nor2_2 _26180_ (.A(_16104_),
    .B(_16106_),
    .Y(_16198_));
 sky130_fd_sc_hd__or3_2 _26181_ (.A(_16196_),
    .B(_16197_),
    .C(_16198_),
    .X(_16199_));
 sky130_fd_sc_hd__o21ai_2 _26182_ (.A1(_16196_),
    .A2(_16197_),
    .B1(_16198_),
    .Y(_16200_));
 sky130_fd_sc_hd__nand3_2 _26183_ (.A(_16178_),
    .B(_16199_),
    .C(_16200_),
    .Y(_16202_));
 sky130_fd_sc_hd__a21o_2 _26184_ (.A1(_16199_),
    .A2(_16200_),
    .B1(_16178_),
    .X(_16203_));
 sky130_fd_sc_hd__and3_2 _26185_ (.A(_16069_),
    .B(_16202_),
    .C(_16203_),
    .X(_16204_));
 sky130_fd_sc_hd__a21oi_2 _26186_ (.A1(_16202_),
    .A2(_16203_),
    .B1(_16069_),
    .Y(_16205_));
 sky130_fd_sc_hd__a211oi_2 _26187_ (.A1(_16109_),
    .A2(_16160_),
    .B1(_16204_),
    .C1(_16205_),
    .Y(_16206_));
 sky130_fd_sc_hd__o211a_2 _26188_ (.A1(_16204_),
    .A2(_16205_),
    .B1(_16109_),
    .C1(_16160_),
    .X(_16207_));
 sky130_fd_sc_hd__nor3_2 _26189_ (.A(_16159_),
    .B(_16206_),
    .C(_16207_),
    .Y(_16208_));
 sky130_fd_sc_hd__o21a_2 _26190_ (.A1(_16206_),
    .A2(_16207_),
    .B1(_16159_),
    .X(_16209_));
 sky130_fd_sc_hd__or3_2 _26191_ (.A(_16118_),
    .B(_16208_),
    .C(_16209_),
    .X(_16210_));
 sky130_fd_sc_hd__o21ai_2 _26192_ (.A1(_16208_),
    .A2(_16209_),
    .B1(_16118_),
    .Y(_16211_));
 sky130_fd_sc_hd__o211ai_2 _26193_ (.A1(_16141_),
    .A2(_16116_),
    .B1(_16210_),
    .C1(_16211_),
    .Y(_16213_));
 sky130_fd_sc_hd__a211o_2 _26194_ (.A1(_16210_),
    .A2(_16211_),
    .B1(_16141_),
    .C1(_16116_),
    .X(_16214_));
 sky130_fd_sc_hd__and2_2 _26195_ (.A(_16213_),
    .B(_16214_),
    .X(_16215_));
 sky130_fd_sc_hd__nor2_2 _26196_ (.A(_16120_),
    .B(_16122_),
    .Y(_16216_));
 sky130_fd_sc_hd__xnor2_2 _26197_ (.A(_16215_),
    .B(_16216_),
    .Y(_16217_));
 sky130_fd_sc_hd__and2b_2 _26198_ (.A_N(_16140_),
    .B(_16217_),
    .X(_16218_));
 sky130_fd_sc_hd__and2b_2 _26199_ (.A_N(_16217_),
    .B(_16140_),
    .X(_16219_));
 sky130_fd_sc_hd__nor2_2 _26200_ (.A(_16218_),
    .B(_16219_),
    .Y(_16220_));
 sky130_fd_sc_hd__nor2_2 _26201_ (.A(_16124_),
    .B(_16127_),
    .Y(_16221_));
 sky130_fd_sc_hd__xnor2_2 _26202_ (.A(_16220_),
    .B(_16221_),
    .Y(_16222_));
 sky130_fd_sc_hd__a21oi_2 _26203_ (.A1(_15570_),
    .A2(_16129_),
    .B1(_16131_),
    .Y(_16224_));
 sky130_fd_sc_hd__o31a_2 _26204_ (.A1(_15573_),
    .A2(_16130_),
    .A3(_16131_),
    .B1(_16224_),
    .X(_16225_));
 sky130_fd_sc_hd__xnor2_2 _26205_ (.A(_16222_),
    .B(_16225_),
    .Y(_16226_));
 sky130_fd_sc_hd__nand2_2 _26206_ (.A(_15823_),
    .B(_15926_),
    .Y(_16227_));
 sky130_fd_sc_hd__nor2_2 _26207_ (.A(_15924_),
    .B(_15925_),
    .Y(_16228_));
 sky130_fd_sc_hd__a31o_2 _26208_ (.A1(_15824_),
    .A2(_15604_),
    .A3(_15850_),
    .B1(_15849_),
    .X(_16229_));
 sky130_fd_sc_hd__nand2_2 _26209_ (.A(_15846_),
    .B(_15845_),
    .Y(_16230_));
 sky130_fd_sc_hd__or3b_2 _26210_ (.A(_15855_),
    .B(_15872_),
    .C_N(_15874_),
    .X(_16231_));
 sky130_fd_sc_hd__and2b_2 _26211_ (.A_N(_15872_),
    .B(_16231_),
    .X(_16232_));
 sky130_fd_sc_hd__a21o_2 _26212_ (.A1(_15836_),
    .A2(_15841_),
    .B1(_15838_),
    .X(_16233_));
 sky130_fd_sc_hd__o2bb2a_2 _26213_ (.A1_N(_15859_),
    .A2_N(_15861_),
    .B1(_15614_),
    .B2(_15858_),
    .X(_16235_));
 sky130_fd_sc_hd__nor2_2 _26214_ (.A(_11570_),
    .B(_15834_),
    .Y(_16236_));
 sky130_fd_sc_hd__buf_1 _26215_ (.A(_15153_),
    .X(_16237_));
 sky130_fd_sc_hd__or3b_2 _26216_ (.A(_15167_),
    .B(_16237_),
    .C_N(_15837_),
    .X(_16238_));
 sky130_fd_sc_hd__a21o_2 _26217_ (.A1(_14388_),
    .A2(_15585_),
    .B1(_15837_),
    .X(_16239_));
 sky130_fd_sc_hd__nand3_2 _26218_ (.A(_16236_),
    .B(_16238_),
    .C(_16239_),
    .Y(_16240_));
 sky130_fd_sc_hd__a21o_2 _26219_ (.A1(_16238_),
    .A2(_16239_),
    .B1(_16236_),
    .X(_16241_));
 sky130_fd_sc_hd__and3b_2 _26220_ (.A_N(_16235_),
    .B(_16240_),
    .C(_16241_),
    .X(_16242_));
 sky130_fd_sc_hd__a21boi_2 _26221_ (.A1(_16240_),
    .A2(_16241_),
    .B1_N(_16235_),
    .Y(_16243_));
 sky130_fd_sc_hd__nor2_2 _26222_ (.A(_16242_),
    .B(_16243_),
    .Y(_16244_));
 sky130_fd_sc_hd__xnor2_2 _26223_ (.A(_16233_),
    .B(_16244_),
    .Y(_16246_));
 sky130_fd_sc_hd__o21bai_2 _26224_ (.A1(_15601_),
    .A2(_15844_),
    .B1_N(_15843_),
    .Y(_16247_));
 sky130_fd_sc_hd__xor2_2 _26225_ (.A(_16246_),
    .B(_16247_),
    .X(_16248_));
 sky130_fd_sc_hd__and2_4 _26226_ (.A(iY[18]),
    .B(iY[50]),
    .X(_16249_));
 sky130_fd_sc_hd__nor2_2 _26227_ (.A(iY[18]),
    .B(iY[50]),
    .Y(_16250_));
 sky130_fd_sc_hd__nor2_2 _26228_ (.A(_16249_),
    .B(_16250_),
    .Y(_16251_));
 sky130_fd_sc_hd__and2_2 _26229_ (.A(iY[17]),
    .B(iY[49]),
    .X(_16252_));
 sky130_fd_sc_hd__o21a_2 _26230_ (.A1(_15593_),
    .A2(_16252_),
    .B1(_15830_),
    .X(_16253_));
 sky130_fd_sc_hd__a31o_2 _26231_ (.A1(_15592_),
    .A2(_15595_),
    .A3(_15830_),
    .B1(_16253_),
    .X(_16254_));
 sky130_fd_sc_hd__xnor2_2 _26232_ (.A(_16251_),
    .B(_16254_),
    .Y(_16255_));
 sky130_fd_sc_hd__buf_1 _26233_ (.A(_16255_),
    .X(_16257_));
 sky130_fd_sc_hd__buf_1 _26234_ (.A(_16257_),
    .X(_16258_));
 sky130_fd_sc_hd__nor2_2 _26235_ (.A(_11578_),
    .B(_16258_),
    .Y(_16259_));
 sky130_fd_sc_hd__xor2_2 _26236_ (.A(_16248_),
    .B(_16259_),
    .X(_16260_));
 sky130_fd_sc_hd__xnor2_2 _26237_ (.A(_16232_),
    .B(_16260_),
    .Y(_16261_));
 sky130_fd_sc_hd__xnor2_2 _26238_ (.A(_16230_),
    .B(_16261_),
    .Y(_16262_));
 sky130_fd_sc_hd__or2_2 _26239_ (.A(_15863_),
    .B(_15870_),
    .X(_16263_));
 sky130_fd_sc_hd__o21ai_2 _26240_ (.A1(_15868_),
    .A2(_15869_),
    .B1(_16263_),
    .Y(_16264_));
 sky130_fd_sc_hd__and2b_2 _26241_ (.A_N(_15885_),
    .B(_15877_),
    .X(_16265_));
 sky130_fd_sc_hd__nor2_2 _26242_ (.A(_15882_),
    .B(_16265_),
    .Y(_16266_));
 sky130_fd_sc_hd__buf_1 _26243_ (.A(_12816_),
    .X(_16268_));
 sky130_fd_sc_hd__nand2_2 _26244_ (.A(_16268_),
    .B(_14411_),
    .Y(_16269_));
 sky130_fd_sc_hd__xor2_2 _26245_ (.A(_15858_),
    .B(_16269_),
    .X(_16270_));
 sky130_fd_sc_hd__buf_6 _26246_ (.A(_14346_),
    .X(_16271_));
 sky130_fd_sc_hd__nor2_2 _26247_ (.A(_16271_),
    .B(_14949_),
    .Y(_16272_));
 sky130_fd_sc_hd__xnor2_2 _26248_ (.A(_16270_),
    .B(_16272_),
    .Y(_16273_));
 sky130_fd_sc_hd__nand2_2 _26249_ (.A(_13244_),
    .B(_13888_),
    .Y(_16274_));
 sky130_fd_sc_hd__nand2_2 _26250_ (.A(_14648_),
    .B(_13543_),
    .Y(_16275_));
 sky130_fd_sc_hd__xnor2_2 _26251_ (.A(_16274_),
    .B(_16275_),
    .Y(_16276_));
 sky130_fd_sc_hd__buf_1 _26252_ (.A(_13501_),
    .X(_16277_));
 sky130_fd_sc_hd__nand2_2 _26253_ (.A(_16277_),
    .B(_14392_),
    .Y(_16279_));
 sky130_fd_sc_hd__xnor2_2 _26254_ (.A(_16276_),
    .B(_16279_),
    .Y(_16280_));
 sky130_fd_sc_hd__o21a_2 _26255_ (.A1(_15866_),
    .A2(_15867_),
    .B1(_15864_),
    .X(_16281_));
 sky130_fd_sc_hd__nor2_2 _26256_ (.A(_16280_),
    .B(_16281_),
    .Y(_16282_));
 sky130_fd_sc_hd__nand2_2 _26257_ (.A(_16280_),
    .B(_16281_),
    .Y(_16283_));
 sky130_fd_sc_hd__or2b_2 _26258_ (.A(_16282_),
    .B_N(_16283_),
    .X(_16284_));
 sky130_fd_sc_hd__xor2_2 _26259_ (.A(_16273_),
    .B(_16284_),
    .X(_16285_));
 sky130_fd_sc_hd__xnor2_2 _26260_ (.A(_16266_),
    .B(_16285_),
    .Y(_16286_));
 sky130_fd_sc_hd__xor2_2 _26261_ (.A(_16264_),
    .B(_16286_),
    .X(_16287_));
 sky130_fd_sc_hd__buf_1 _26262_ (.A(_14983_),
    .X(_16288_));
 sky130_fd_sc_hd__or3b_2 _26263_ (.A(_12852_),
    .B(_15647_),
    .C_N(_15637_),
    .X(_16290_));
 sky130_fd_sc_hd__o31ai_2 _26264_ (.A1(_14626_),
    .A2(_16288_),
    .A3(_15878_),
    .B1(_16290_),
    .Y(_16291_));
 sky130_fd_sc_hd__buf_1 _26265_ (.A(_14999_),
    .X(_16292_));
 sky130_fd_sc_hd__and3_2 _26266_ (.A(_14980_),
    .B(_16292_),
    .C(_15891_),
    .X(_16293_));
 sky130_fd_sc_hd__a31o_2 _26267_ (.A1(_15887_),
    .A2(_15208_),
    .A3(_15892_),
    .B1(_16293_),
    .X(_16294_));
 sky130_fd_sc_hd__or4_2 _26268_ (.A(_12773_),
    .B(_12850_),
    .C(_13934_),
    .D(_14987_),
    .X(_16295_));
 sky130_fd_sc_hd__a22o_2 _26269_ (.A1(_12846_),
    .A2(_13938_),
    .B1(_15208_),
    .B2(_14634_),
    .X(_16296_));
 sky130_fd_sc_hd__nand2_2 _26270_ (.A(_16295_),
    .B(_16296_),
    .Y(_16297_));
 sky130_fd_sc_hd__nor2_2 _26271_ (.A(_14625_),
    .B(_15211_),
    .Y(_16298_));
 sky130_fd_sc_hd__xnor2_2 _26272_ (.A(_16297_),
    .B(_16298_),
    .Y(_16299_));
 sky130_fd_sc_hd__xor2_2 _26273_ (.A(_16294_),
    .B(_16299_),
    .X(_16301_));
 sky130_fd_sc_hd__and2_2 _26274_ (.A(_16291_),
    .B(_16301_),
    .X(_16302_));
 sky130_fd_sc_hd__nor2_2 _26275_ (.A(_16291_),
    .B(_16301_),
    .Y(_16303_));
 sky130_fd_sc_hd__nor2_2 _26276_ (.A(_16302_),
    .B(_16303_),
    .Y(_16304_));
 sky130_fd_sc_hd__nor2_2 _26277_ (.A(_14356_),
    .B(_15005_),
    .Y(_16305_));
 sky130_fd_sc_hd__or4b_2 _26278_ (.A(_12248_),
    .B(_15219_),
    .C(_15220_),
    .D_N(_15891_),
    .X(_16306_));
 sky130_fd_sc_hd__a32o_2 _26279_ (.A1(_14649_),
    .A2(_15224_),
    .A3(_15226_),
    .B1(_14980_),
    .B2(_15679_),
    .X(_16307_));
 sky130_fd_sc_hd__nand3_2 _26280_ (.A(_16305_),
    .B(_16306_),
    .C(_16307_),
    .Y(_16308_));
 sky130_fd_sc_hd__a21o_2 _26281_ (.A1(_16306_),
    .A2(_16307_),
    .B1(_16305_),
    .X(_16309_));
 sky130_fd_sc_hd__and2_2 _26282_ (.A(_16308_),
    .B(_16309_),
    .X(_16310_));
 sky130_fd_sc_hd__buf_1 _26283_ (.A(_15668_),
    .X(_16312_));
 sky130_fd_sc_hd__nor2_2 _26284_ (.A(_11791_),
    .B(_16312_),
    .Y(_16313_));
 sky130_fd_sc_hd__nand2_2 _26285_ (.A(_11583_),
    .B(_15899_),
    .Y(_16314_));
 sky130_fd_sc_hd__or2b_2 _26286_ (.A(_15664_),
    .B_N(_15896_),
    .X(_16315_));
 sky130_fd_sc_hd__a21o_2 _26287_ (.A1(_15663_),
    .A2(_15667_),
    .B1(_16315_),
    .X(_16316_));
 sky130_fd_sc_hd__xnor2_2 _26288_ (.A(iX[18]),
    .B(iX[50]),
    .Y(_16317_));
 sky130_fd_sc_hd__and2b_2 _26289_ (.A_N(_16317_),
    .B(_15894_),
    .X(_16318_));
 sky130_fd_sc_hd__nand2_2 _26290_ (.A(_16316_),
    .B(_16318_),
    .Y(_16319_));
 sky130_fd_sc_hd__a21bo_2 _26291_ (.A1(_15894_),
    .A2(_16316_),
    .B1_N(_16317_),
    .X(_16320_));
 sky130_fd_sc_hd__and3_2 _26292_ (.A(_11379_),
    .B(_16319_),
    .C(_16320_),
    .X(_16321_));
 sky130_fd_sc_hd__xnor2_2 _26293_ (.A(_16314_),
    .B(_16321_),
    .Y(_16323_));
 sky130_fd_sc_hd__xor2_2 _26294_ (.A(_16313_),
    .B(_16323_),
    .X(_16324_));
 sky130_fd_sc_hd__o21a_2 _26295_ (.A1(_15901_),
    .A2(_15904_),
    .B1(_16324_),
    .X(_16325_));
 sky130_fd_sc_hd__or3_2 _26296_ (.A(_15901_),
    .B(_15904_),
    .C(_16324_),
    .X(_16326_));
 sky130_fd_sc_hd__and2b_2 _26297_ (.A_N(_16325_),
    .B(_16326_),
    .X(_16327_));
 sky130_fd_sc_hd__xnor2_2 _26298_ (.A(_16310_),
    .B(_16327_),
    .Y(_16328_));
 sky130_fd_sc_hd__and2_2 _26299_ (.A(_15907_),
    .B(_15908_),
    .X(_16329_));
 sky130_fd_sc_hd__a21oi_2 _26300_ (.A1(_15893_),
    .A2(_15909_),
    .B1(_16329_),
    .Y(_16330_));
 sky130_fd_sc_hd__xnor2_2 _26301_ (.A(_16328_),
    .B(_16330_),
    .Y(_16331_));
 sky130_fd_sc_hd__xnor2_2 _26302_ (.A(_16304_),
    .B(_16331_),
    .Y(_16332_));
 sky130_fd_sc_hd__nor2_2 _26303_ (.A(_15910_),
    .B(_15911_),
    .Y(_16334_));
 sky130_fd_sc_hd__a21o_2 _26304_ (.A1(_15886_),
    .A2(_15912_),
    .B1(_16334_),
    .X(_16335_));
 sky130_fd_sc_hd__xor2_2 _26305_ (.A(_16332_),
    .B(_16335_),
    .X(_16336_));
 sky130_fd_sc_hd__xor2_2 _26306_ (.A(_16287_),
    .B(_16336_),
    .X(_16337_));
 sky130_fd_sc_hd__and2b_2 _26307_ (.A_N(_15913_),
    .B(_15914_),
    .X(_16338_));
 sky130_fd_sc_hd__a21oi_2 _26308_ (.A1(_15876_),
    .A2(_15915_),
    .B1(_16338_),
    .Y(_16339_));
 sky130_fd_sc_hd__xnor2_2 _26309_ (.A(_16337_),
    .B(_16339_),
    .Y(_16340_));
 sky130_fd_sc_hd__xnor2_2 _26310_ (.A(_16262_),
    .B(_16340_),
    .Y(_16341_));
 sky130_fd_sc_hd__and2b_2 _26311_ (.A_N(_15919_),
    .B(_15916_),
    .X(_16342_));
 sky130_fd_sc_hd__a21oi_2 _26312_ (.A1(_15853_),
    .A2(_15920_),
    .B1(_16342_),
    .Y(_16343_));
 sky130_fd_sc_hd__xor2_2 _26313_ (.A(_16341_),
    .B(_16343_),
    .X(_16345_));
 sky130_fd_sc_hd__xnor2_2 _26314_ (.A(_16229_),
    .B(_16345_),
    .Y(_16346_));
 sky130_fd_sc_hd__and2b_2 _26315_ (.A_N(_15921_),
    .B(_15922_),
    .X(_16347_));
 sky130_fd_sc_hd__a21oi_2 _26316_ (.A1(_15606_),
    .A2(_15923_),
    .B1(_16347_),
    .Y(_16348_));
 sky130_fd_sc_hd__xor2_2 _26317_ (.A(_16346_),
    .B(_16348_),
    .X(_16349_));
 sky130_fd_sc_hd__xor2_2 _26318_ (.A(_16228_),
    .B(_16349_),
    .X(_16350_));
 sky130_fd_sc_hd__xnor2_2 _26319_ (.A(_16227_),
    .B(_16350_),
    .Y(_16351_));
 sky130_fd_sc_hd__and3b_2 _26320_ (.A_N(_15708_),
    .B(_15927_),
    .C(_15707_),
    .X(_16352_));
 sky130_fd_sc_hd__a31o_2 _26321_ (.A1(_15579_),
    .A2(_15710_),
    .A3(_15927_),
    .B1(_16352_),
    .X(_16353_));
 sky130_fd_sc_hd__xnor2_2 _26322_ (.A(_16351_),
    .B(_16353_),
    .Y(_16354_));
 sky130_fd_sc_hd__or3_2 _26323_ (.A(_16019_),
    .B(_16020_),
    .C(_16022_),
    .X(_16356_));
 sky130_fd_sc_hd__inv_2 _26324_ (.A(_16019_),
    .Y(_16357_));
 sky130_fd_sc_hd__inv_2 _26325_ (.A(_15995_),
    .Y(_16358_));
 sky130_fd_sc_hd__or2b_2 _26326_ (.A(_15941_),
    .B_N(_15940_),
    .X(_16359_));
 sky130_fd_sc_hd__nand2_2 _26327_ (.A(_15942_),
    .B(_15947_),
    .Y(_16360_));
 sky130_fd_sc_hd__and4_2 _26328_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[47]),
    .D(iX[48]),
    .X(_16361_));
 sky130_fd_sc_hd__a22oi_2 _26329_ (.A1(iY[35]),
    .A2(iX[47]),
    .B1(iX[48]),
    .B2(iY[34]),
    .Y(_16362_));
 sky130_fd_sc_hd__nor2_2 _26330_ (.A(_16361_),
    .B(_16362_),
    .Y(_16363_));
 sky130_fd_sc_hd__nand2_2 _26331_ (.A(iY[33]),
    .B(iX[49]),
    .Y(_16364_));
 sky130_fd_sc_hd__xnor2_2 _26332_ (.A(_16363_),
    .B(_16364_),
    .Y(_16365_));
 sky130_fd_sc_hd__o21ba_2 _26333_ (.A1(_15936_),
    .A2(_15938_),
    .B1_N(_15935_),
    .X(_16367_));
 sky130_fd_sc_hd__xnor2_2 _26334_ (.A(_16365_),
    .B(_16367_),
    .Y(_16368_));
 sky130_fd_sc_hd__and4_2 _26335_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[46]),
    .D(iX[50]),
    .X(_16369_));
 sky130_fd_sc_hd__a22oi_2 _26336_ (.A1(iY[36]),
    .A2(iX[46]),
    .B1(iX[50]),
    .B2(iY[32]),
    .Y(_16370_));
 sky130_fd_sc_hd__nor2_2 _26337_ (.A(_16369_),
    .B(_16370_),
    .Y(_16371_));
 sky130_fd_sc_hd__nand2_2 _26338_ (.A(iY[37]),
    .B(iX[45]),
    .Y(_16372_));
 sky130_fd_sc_hd__xnor2_2 _26339_ (.A(_16371_),
    .B(_16372_),
    .Y(_16373_));
 sky130_fd_sc_hd__xnor2_2 _26340_ (.A(_16368_),
    .B(_16373_),
    .Y(_16374_));
 sky130_fd_sc_hd__a21o_2 _26341_ (.A1(_16359_),
    .A2(_16360_),
    .B1(_16374_),
    .X(_16375_));
 sky130_fd_sc_hd__nand3_2 _26342_ (.A(_16359_),
    .B(_16360_),
    .C(_16374_),
    .Y(_16376_));
 sky130_fd_sc_hd__o21ba_2 _26343_ (.A1(_15955_),
    .A2(_15957_),
    .B1_N(_15954_),
    .X(_16378_));
 sky130_fd_sc_hd__o21ba_2 _26344_ (.A1(_15944_),
    .A2(_15946_),
    .B1_N(_15943_),
    .X(_16379_));
 sky130_fd_sc_hd__and4_2 _26345_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[43]),
    .D(iX[44]),
    .X(_16380_));
 sky130_fd_sc_hd__a22oi_2 _26346_ (.A1(iY[39]),
    .A2(iX[43]),
    .B1(iX[44]),
    .B2(iY[38]),
    .Y(_16381_));
 sky130_fd_sc_hd__nor2_2 _26347_ (.A(_16380_),
    .B(_16381_),
    .Y(_16382_));
 sky130_fd_sc_hd__nand2_2 _26348_ (.A(iY[40]),
    .B(iX[42]),
    .Y(_16383_));
 sky130_fd_sc_hd__xnor2_2 _26349_ (.A(_16382_),
    .B(_16383_),
    .Y(_16384_));
 sky130_fd_sc_hd__xnor2_2 _26350_ (.A(_16379_),
    .B(_16384_),
    .Y(_16385_));
 sky130_fd_sc_hd__xnor2_2 _26351_ (.A(_16378_),
    .B(_16385_),
    .Y(_16386_));
 sky130_fd_sc_hd__nand3_2 _26352_ (.A(_16375_),
    .B(_16376_),
    .C(_16386_),
    .Y(_16387_));
 sky130_fd_sc_hd__a21o_2 _26353_ (.A1(_16375_),
    .A2(_16376_),
    .B1(_16386_),
    .X(_16389_));
 sky130_fd_sc_hd__nand2_2 _26354_ (.A(_16387_),
    .B(_16389_),
    .Y(_16390_));
 sky130_fd_sc_hd__nand2_2 _26355_ (.A(_15949_),
    .B(_15962_),
    .Y(_16391_));
 sky130_fd_sc_hd__xnor2_2 _26356_ (.A(_16390_),
    .B(_16391_),
    .Y(_16392_));
 sky130_fd_sc_hd__and2b_2 _26357_ (.A_N(_15982_),
    .B(_15981_),
    .X(_16393_));
 sky130_fd_sc_hd__or2b_2 _26358_ (.A(_15953_),
    .B_N(_15958_),
    .X(_16394_));
 sky130_fd_sc_hd__or2b_2 _26359_ (.A(_15952_),
    .B_N(_15959_),
    .X(_16395_));
 sky130_fd_sc_hd__and4_2 _26360_ (.A(iX[37]),
    .B(iX[38]),
    .C(iY[44]),
    .D(iY[45]),
    .X(_16396_));
 sky130_fd_sc_hd__a22oi_2 _26361_ (.A1(iX[38]),
    .A2(iY[44]),
    .B1(iY[45]),
    .B2(iX[37]),
    .Y(_16397_));
 sky130_fd_sc_hd__nor2_2 _26362_ (.A(_16396_),
    .B(_16397_),
    .Y(_16398_));
 sky130_fd_sc_hd__nand2_2 _26363_ (.A(iX[36]),
    .B(iY[46]),
    .Y(_16400_));
 sky130_fd_sc_hd__xnor2_2 _26364_ (.A(_16398_),
    .B(_16400_),
    .Y(_16401_));
 sky130_fd_sc_hd__and4_2 _26365_ (.A(iX[40]),
    .B(iX[41]),
    .C(iY[41]),
    .D(iY[42]),
    .X(_16402_));
 sky130_fd_sc_hd__a22oi_2 _26366_ (.A1(iX[41]),
    .A2(iY[41]),
    .B1(iY[42]),
    .B2(iX[40]),
    .Y(_16403_));
 sky130_fd_sc_hd__nor2_2 _26367_ (.A(_16402_),
    .B(_16403_),
    .Y(_16404_));
 sky130_fd_sc_hd__nand2_2 _26368_ (.A(iX[39]),
    .B(iY[43]),
    .Y(_16405_));
 sky130_fd_sc_hd__xnor2_2 _26369_ (.A(_16404_),
    .B(_16405_),
    .Y(_16406_));
 sky130_fd_sc_hd__o21ba_2 _26370_ (.A1(_15978_),
    .A2(_15980_),
    .B1_N(_15977_),
    .X(_16407_));
 sky130_fd_sc_hd__xnor2_2 _26371_ (.A(_16406_),
    .B(_16407_),
    .Y(_16408_));
 sky130_fd_sc_hd__xnor2_2 _26372_ (.A(_16401_),
    .B(_16408_),
    .Y(_16409_));
 sky130_fd_sc_hd__a21o_2 _26373_ (.A1(_16394_),
    .A2(_16395_),
    .B1(_16409_),
    .X(_16411_));
 sky130_fd_sc_hd__nand3_2 _26374_ (.A(_16394_),
    .B(_16395_),
    .C(_16409_),
    .Y(_16412_));
 sky130_fd_sc_hd__o211ai_2 _26375_ (.A1(_16393_),
    .A2(_15985_),
    .B1(_16411_),
    .C1(_16412_),
    .Y(_16413_));
 sky130_fd_sc_hd__a211o_2 _26376_ (.A1(_16411_),
    .A2(_16412_),
    .B1(_16393_),
    .C1(_15985_),
    .X(_16414_));
 sky130_fd_sc_hd__and3_2 _26377_ (.A(_16392_),
    .B(_16413_),
    .C(_16414_),
    .X(_16415_));
 sky130_fd_sc_hd__inv_2 _26378_ (.A(_16415_),
    .Y(_16416_));
 sky130_fd_sc_hd__a21o_2 _26379_ (.A1(_16413_),
    .A2(_16414_),
    .B1(_16392_),
    .X(_16417_));
 sky130_fd_sc_hd__o211a_2 _26380_ (.A1(_15965_),
    .A2(_15992_),
    .B1(_16416_),
    .C1(_16417_),
    .X(_16418_));
 sky130_fd_sc_hd__a211oi_2 _26381_ (.A1(_16416_),
    .A2(_16417_),
    .B1(_15965_),
    .C1(_15992_),
    .Y(_16419_));
 sky130_fd_sc_hd__and2_2 _26382_ (.A(_16007_),
    .B(_16004_),
    .X(_16420_));
 sky130_fd_sc_hd__o21ba_2 _26383_ (.A1(_15973_),
    .A2(_15975_),
    .B1_N(_15971_),
    .X(_16422_));
 sky130_fd_sc_hd__and4_2 _26384_ (.A(iX[34]),
    .B(iX[35]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_16423_));
 sky130_fd_sc_hd__a22oi_2 _26385_ (.A1(iX[35]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[34]),
    .Y(_16424_));
 sky130_fd_sc_hd__nor2_2 _26386_ (.A(_16423_),
    .B(_16424_),
    .Y(_16425_));
 sky130_fd_sc_hd__nand2_2 _26387_ (.A(iX[33]),
    .B(iY[49]),
    .Y(_16426_));
 sky130_fd_sc_hd__xnor2_2 _26388_ (.A(_16425_),
    .B(_16426_),
    .Y(_16427_));
 sky130_fd_sc_hd__xnor2_2 _26389_ (.A(_16422_),
    .B(_16427_),
    .Y(_16428_));
 sky130_fd_sc_hd__a31oi_2 _26390_ (.A1(iX[32]),
    .A2(iY[49]),
    .A3(_15999_),
    .B1(_15998_),
    .Y(_16429_));
 sky130_fd_sc_hd__or2b_2 _26391_ (.A(_16428_),
    .B_N(_16429_),
    .X(_16430_));
 sky130_fd_sc_hd__or2b_2 _26392_ (.A(_16429_),
    .B_N(_16428_),
    .X(_16431_));
 sky130_fd_sc_hd__nand2_2 _26393_ (.A(_16430_),
    .B(_16431_),
    .Y(_16433_));
 sky130_fd_sc_hd__a21oi_2 _26394_ (.A1(_16006_),
    .A2(_16004_),
    .B1(_16003_),
    .Y(_16434_));
 sky130_fd_sc_hd__xor2_2 _26395_ (.A(_16433_),
    .B(_16434_),
    .X(_16435_));
 sky130_fd_sc_hd__and2_2 _26396_ (.A(iX[32]),
    .B(iY[50]),
    .X(_16436_));
 sky130_fd_sc_hd__nor2_2 _26397_ (.A(_16435_),
    .B(_16436_),
    .Y(_16437_));
 sky130_fd_sc_hd__and2_2 _26398_ (.A(_16435_),
    .B(_16436_),
    .X(_16438_));
 sky130_fd_sc_hd__or2_2 _26399_ (.A(_16437_),
    .B(_16438_),
    .X(_16439_));
 sky130_fd_sc_hd__a21oi_2 _26400_ (.A1(_15988_),
    .A2(_15990_),
    .B1(_16439_),
    .Y(_16440_));
 sky130_fd_sc_hd__and3_2 _26401_ (.A(_15988_),
    .B(_15990_),
    .C(_16439_),
    .X(_16441_));
 sky130_fd_sc_hd__nor2_2 _26402_ (.A(_16440_),
    .B(_16441_),
    .Y(_16442_));
 sky130_fd_sc_hd__xnor2_2 _26403_ (.A(_16420_),
    .B(_16442_),
    .Y(_16444_));
 sky130_fd_sc_hd__o21ai_2 _26404_ (.A1(_16418_),
    .A2(_16419_),
    .B1(_16444_),
    .Y(_16445_));
 sky130_fd_sc_hd__or3_2 _26405_ (.A(_16418_),
    .B(_16419_),
    .C(_16444_),
    .X(_16446_));
 sky130_fd_sc_hd__o211a_2 _26406_ (.A1(_16358_),
    .A2(_16015_),
    .B1(_16445_),
    .C1(_16446_),
    .X(_16447_));
 sky130_fd_sc_hd__a211oi_2 _26407_ (.A1(_16445_),
    .A2(_16446_),
    .B1(_16358_),
    .C1(_16015_),
    .Y(_16448_));
 sky130_fd_sc_hd__nor2_2 _26408_ (.A(_16447_),
    .B(_16448_),
    .Y(_16449_));
 sky130_fd_sc_hd__o21a_2 _26409_ (.A1(_15789_),
    .A2(_16012_),
    .B1(_16010_),
    .X(_16450_));
 sky130_fd_sc_hd__xor2_2 _26410_ (.A(_16449_),
    .B(_16450_),
    .X(_16451_));
 sky130_fd_sc_hd__a21oi_2 _26411_ (.A1(_16017_),
    .A2(_16357_),
    .B1(_16451_),
    .Y(_16452_));
 sky130_fd_sc_hd__and3_2 _26412_ (.A(_16017_),
    .B(_16357_),
    .C(_16451_),
    .X(_16453_));
 sky130_fd_sc_hd__nor3_2 _26413_ (.A(_16356_),
    .B(_16452_),
    .C(_16453_),
    .Y(_16455_));
 sky130_fd_sc_hd__o21a_2 _26414_ (.A1(_16452_),
    .A2(_16453_),
    .B1(_16356_),
    .X(_16456_));
 sky130_fd_sc_hd__o21ba_2 _26415_ (.A1(_16455_),
    .A2(_16456_),
    .B1_N(_16024_),
    .X(_16457_));
 sky130_fd_sc_hd__nor3b_2 _26416_ (.A(_16455_),
    .B(_16456_),
    .C_N(_16024_),
    .Y(_16458_));
 sky130_fd_sc_hd__and3_2 _26417_ (.A(_15713_),
    .B(_15806_),
    .C(_16026_),
    .X(_16459_));
 sky130_fd_sc_hd__a21o_2 _26418_ (.A1(_16028_),
    .A2(_16032_),
    .B1(_16029_),
    .X(_16460_));
 sky130_fd_sc_hd__or3_2 _26419_ (.A(_16458_),
    .B(_16459_),
    .C(_16460_),
    .X(_16461_));
 sky130_fd_sc_hd__o22ai_2 _26420_ (.A1(_16458_),
    .A2(_16457_),
    .B1(_16459_),
    .B2(_16460_),
    .Y(_16462_));
 sky130_fd_sc_hd__o21a_2 _26421_ (.A1(_16457_),
    .A2(_16461_),
    .B1(_16462_),
    .X(_16463_));
 sky130_fd_sc_hd__xor2_2 _26422_ (.A(_16354_),
    .B(_16463_),
    .X(_16464_));
 sky130_fd_sc_hd__xor2_2 _26423_ (.A(oO[18]),
    .B(_16464_),
    .X(_16466_));
 sky130_fd_sc_hd__and2b_2 _26424_ (.A_N(_15930_),
    .B(_16034_),
    .X(_16467_));
 sky130_fd_sc_hd__and2b_2 _26425_ (.A_N(oO[17]),
    .B(_16035_),
    .X(_16468_));
 sky130_fd_sc_hd__nor2_2 _26426_ (.A(_16467_),
    .B(_16468_),
    .Y(_16469_));
 sky130_fd_sc_hd__xor2_2 _26427_ (.A(_16466_),
    .B(_16469_),
    .X(_16470_));
 sky130_fd_sc_hd__or2b_2 _26428_ (.A(_16036_),
    .B_N(_16040_),
    .X(_16471_));
 sky130_fd_sc_hd__or3b_2 _26429_ (.A(_15578_),
    .B(_16041_),
    .C_N(_15810_),
    .X(_16472_));
 sky130_fd_sc_hd__a311o_2 _26430_ (.A1(_16037_),
    .A2(_16039_),
    .A3(_16036_),
    .B1(_15814_),
    .C1(_15813_),
    .X(_16473_));
 sky130_fd_sc_hd__and3_2 _26431_ (.A(_16471_),
    .B(_16472_),
    .C(_16473_),
    .X(_16474_));
 sky130_fd_sc_hd__or2_2 _26432_ (.A(_16470_),
    .B(_16474_),
    .X(_16475_));
 sky130_fd_sc_hd__nand2_2 _26433_ (.A(_16470_),
    .B(_16474_),
    .Y(_16477_));
 sky130_fd_sc_hd__and3_2 _26434_ (.A(_16226_),
    .B(_16475_),
    .C(_16477_),
    .X(_16478_));
 sky130_fd_sc_hd__a21oi_2 _26435_ (.A1(_16475_),
    .A2(_16477_),
    .B1(_16226_),
    .Y(_16479_));
 sky130_fd_sc_hd__nor2_2 _26436_ (.A(_16478_),
    .B(_16479_),
    .Y(_16480_));
 sky130_fd_sc_hd__a211o_2 _26437_ (.A1(_15461_),
    .A2(_15466_),
    .B1(_15818_),
    .C1(_16138_),
    .X(_16481_));
 sky130_fd_sc_hd__a21oi_2 _26438_ (.A1(_15816_),
    .A2(_16137_),
    .B1(_16135_),
    .Y(_16482_));
 sky130_fd_sc_hd__nand2_2 _26439_ (.A(_16481_),
    .B(_16482_),
    .Y(_16483_));
 sky130_fd_sc_hd__xor2_2 _26440_ (.A(_16480_),
    .B(_16483_),
    .X(oO[50]));
 sky130_fd_sc_hd__o21a_2 _26441_ (.A1(_16467_),
    .A2(_16468_),
    .B1(_16466_),
    .X(_16484_));
 sky130_fd_sc_hd__and2b_2 _26442_ (.A_N(_16450_),
    .B(_16449_),
    .X(_16485_));
 sky130_fd_sc_hd__and3_2 _26443_ (.A(_16387_),
    .B(_16389_),
    .C(_16391_),
    .X(_16487_));
 sky130_fd_sc_hd__and2b_2 _26444_ (.A_N(_16407_),
    .B(_16406_),
    .X(_16488_));
 sky130_fd_sc_hd__and2_2 _26445_ (.A(_16401_),
    .B(_16408_),
    .X(_16489_));
 sky130_fd_sc_hd__or2b_2 _26446_ (.A(_16379_),
    .B_N(_16384_),
    .X(_16490_));
 sky130_fd_sc_hd__or2b_2 _26447_ (.A(_16378_),
    .B_N(_16385_),
    .X(_16491_));
 sky130_fd_sc_hd__and4_2 _26448_ (.A(iX[38]),
    .B(iX[39]),
    .C(iY[44]),
    .D(iY[45]),
    .X(_16492_));
 sky130_fd_sc_hd__a22oi_2 _26449_ (.A1(iX[39]),
    .A2(iY[44]),
    .B1(iY[45]),
    .B2(iX[38]),
    .Y(_16493_));
 sky130_fd_sc_hd__nor2_2 _26450_ (.A(_16492_),
    .B(_16493_),
    .Y(_16494_));
 sky130_fd_sc_hd__nand2_2 _26451_ (.A(iX[37]),
    .B(iY[46]),
    .Y(_16495_));
 sky130_fd_sc_hd__xnor2_2 _26452_ (.A(_16494_),
    .B(_16495_),
    .Y(_16496_));
 sky130_fd_sc_hd__and4_2 _26453_ (.A(iX[41]),
    .B(iY[41]),
    .C(iX[42]),
    .D(iY[42]),
    .X(_16498_));
 sky130_fd_sc_hd__a22oi_2 _26454_ (.A1(iY[41]),
    .A2(iX[42]),
    .B1(iY[42]),
    .B2(iX[41]),
    .Y(_16499_));
 sky130_fd_sc_hd__nor2_2 _26455_ (.A(_16498_),
    .B(_16499_),
    .Y(_16500_));
 sky130_fd_sc_hd__nand2_2 _26456_ (.A(iX[40]),
    .B(iY[43]),
    .Y(_16501_));
 sky130_fd_sc_hd__xnor2_2 _26457_ (.A(_16500_),
    .B(_16501_),
    .Y(_16502_));
 sky130_fd_sc_hd__o21ba_2 _26458_ (.A1(_16403_),
    .A2(_16405_),
    .B1_N(_16402_),
    .X(_16503_));
 sky130_fd_sc_hd__xnor2_2 _26459_ (.A(_16502_),
    .B(_16503_),
    .Y(_16504_));
 sky130_fd_sc_hd__and2_2 _26460_ (.A(_16496_),
    .B(_16504_),
    .X(_16505_));
 sky130_fd_sc_hd__nor2_2 _26461_ (.A(_16496_),
    .B(_16504_),
    .Y(_16506_));
 sky130_fd_sc_hd__or2_2 _26462_ (.A(_16505_),
    .B(_16506_),
    .X(_16507_));
 sky130_fd_sc_hd__a21o_2 _26463_ (.A1(_16490_),
    .A2(_16491_),
    .B1(_16507_),
    .X(_16509_));
 sky130_fd_sc_hd__nand3_2 _26464_ (.A(_16490_),
    .B(_16491_),
    .C(_16507_),
    .Y(_16510_));
 sky130_fd_sc_hd__o211ai_2 _26465_ (.A1(_16488_),
    .A2(_16489_),
    .B1(_16509_),
    .C1(_16510_),
    .Y(_16511_));
 sky130_fd_sc_hd__a211o_2 _26466_ (.A1(_16509_),
    .A2(_16510_),
    .B1(_16488_),
    .C1(_16489_),
    .X(_16512_));
 sky130_fd_sc_hd__or2b_2 _26467_ (.A(_16367_),
    .B_N(_16365_),
    .X(_16513_));
 sky130_fd_sc_hd__nand2_2 _26468_ (.A(_16368_),
    .B(_16373_),
    .Y(_16514_));
 sky130_fd_sc_hd__and4_2 _26469_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[48]),
    .D(iX[49]),
    .X(_16515_));
 sky130_fd_sc_hd__a22oi_2 _26470_ (.A1(iY[35]),
    .A2(iX[48]),
    .B1(iX[49]),
    .B2(iY[34]),
    .Y(_16516_));
 sky130_fd_sc_hd__nor2_2 _26471_ (.A(_16515_),
    .B(_16516_),
    .Y(_16517_));
 sky130_fd_sc_hd__nand2_2 _26472_ (.A(iY[33]),
    .B(iX[50]),
    .Y(_16518_));
 sky130_fd_sc_hd__xnor2_2 _26473_ (.A(_16517_),
    .B(_16518_),
    .Y(_16520_));
 sky130_fd_sc_hd__o21ba_2 _26474_ (.A1(_16362_),
    .A2(_16364_),
    .B1_N(_16361_),
    .X(_16521_));
 sky130_fd_sc_hd__xnor2_2 _26475_ (.A(_16520_),
    .B(_16521_),
    .Y(_16522_));
 sky130_fd_sc_hd__and4_2 _26476_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[47]),
    .D(iX[51]),
    .X(_16523_));
 sky130_fd_sc_hd__a22oi_2 _26477_ (.A1(iY[36]),
    .A2(iX[47]),
    .B1(iX[51]),
    .B2(iY[32]),
    .Y(_16524_));
 sky130_fd_sc_hd__nor2_2 _26478_ (.A(_16523_),
    .B(_16524_),
    .Y(_16525_));
 sky130_fd_sc_hd__nand2_2 _26479_ (.A(iY[37]),
    .B(iX[46]),
    .Y(_16526_));
 sky130_fd_sc_hd__xnor2_2 _26480_ (.A(_16525_),
    .B(_16526_),
    .Y(_16527_));
 sky130_fd_sc_hd__xnor2_2 _26481_ (.A(_16522_),
    .B(_16527_),
    .Y(_16528_));
 sky130_fd_sc_hd__a21o_2 _26482_ (.A1(_16513_),
    .A2(_16514_),
    .B1(_16528_),
    .X(_16529_));
 sky130_fd_sc_hd__nand3_2 _26483_ (.A(_16513_),
    .B(_16514_),
    .C(_16528_),
    .Y(_16531_));
 sky130_fd_sc_hd__o21ba_2 _26484_ (.A1(_16381_),
    .A2(_16383_),
    .B1_N(_16380_),
    .X(_16532_));
 sky130_fd_sc_hd__o21ba_2 _26485_ (.A1(_16370_),
    .A2(_16372_),
    .B1_N(_16369_),
    .X(_16533_));
 sky130_fd_sc_hd__and4_2 _26486_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[44]),
    .D(iX[45]),
    .X(_16534_));
 sky130_fd_sc_hd__a22oi_2 _26487_ (.A1(iY[39]),
    .A2(iX[44]),
    .B1(iX[45]),
    .B2(iY[38]),
    .Y(_16535_));
 sky130_fd_sc_hd__nor2_2 _26488_ (.A(_16534_),
    .B(_16535_),
    .Y(_16536_));
 sky130_fd_sc_hd__nand2_2 _26489_ (.A(iY[40]),
    .B(iX[43]),
    .Y(_16537_));
 sky130_fd_sc_hd__xnor2_2 _26490_ (.A(_16536_),
    .B(_16537_),
    .Y(_16538_));
 sky130_fd_sc_hd__xnor2_2 _26491_ (.A(_16533_),
    .B(_16538_),
    .Y(_16539_));
 sky130_fd_sc_hd__xnor2_2 _26492_ (.A(_16532_),
    .B(_16539_),
    .Y(_16540_));
 sky130_fd_sc_hd__nand3_2 _26493_ (.A(_16529_),
    .B(_16531_),
    .C(_16540_),
    .Y(_16542_));
 sky130_fd_sc_hd__a21o_2 _26494_ (.A1(_16529_),
    .A2(_16531_),
    .B1(_16540_),
    .X(_16543_));
 sky130_fd_sc_hd__nand2_2 _26495_ (.A(_16542_),
    .B(_16543_),
    .Y(_16544_));
 sky130_fd_sc_hd__nand2_2 _26496_ (.A(_16375_),
    .B(_16387_),
    .Y(_16545_));
 sky130_fd_sc_hd__xnor2_2 _26497_ (.A(_16544_),
    .B(_16545_),
    .Y(_16546_));
 sky130_fd_sc_hd__a21o_2 _26498_ (.A1(_16511_),
    .A2(_16512_),
    .B1(_16546_),
    .X(_16547_));
 sky130_fd_sc_hd__and3_2 _26499_ (.A(_16546_),
    .B(_16511_),
    .C(_16512_),
    .X(_16548_));
 sky130_fd_sc_hd__inv_2 _26500_ (.A(_16548_),
    .Y(_16549_));
 sky130_fd_sc_hd__o211ai_2 _26501_ (.A1(_16487_),
    .A2(_16415_),
    .B1(_16547_),
    .C1(_16549_),
    .Y(_16550_));
 sky130_fd_sc_hd__a211o_2 _26502_ (.A1(_16547_),
    .A2(_16549_),
    .B1(_16487_),
    .C1(_16415_),
    .X(_16551_));
 sky130_fd_sc_hd__nand2_2 _26503_ (.A(_16550_),
    .B(_16551_),
    .Y(_16553_));
 sky130_fd_sc_hd__nor2_2 _26504_ (.A(_16433_),
    .B(_16434_),
    .Y(_16554_));
 sky130_fd_sc_hd__nand2_2 _26505_ (.A(_16411_),
    .B(_16413_),
    .Y(_16555_));
 sky130_fd_sc_hd__a22oi_2 _26506_ (.A1(iX[33]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[32]),
    .Y(_16556_));
 sky130_fd_sc_hd__and3_2 _26507_ (.A(iX[33]),
    .B(iY[51]),
    .C(_16436_),
    .X(_16557_));
 sky130_fd_sc_hd__or2b_2 _26508_ (.A(_16422_),
    .B_N(_16427_),
    .X(_16558_));
 sky130_fd_sc_hd__a31o_2 _26509_ (.A1(iX[33]),
    .A2(iY[49]),
    .A3(_16425_),
    .B1(_16423_),
    .X(_16559_));
 sky130_fd_sc_hd__o21ba_2 _26510_ (.A1(_16397_),
    .A2(_16400_),
    .B1_N(_16396_),
    .X(_16560_));
 sky130_fd_sc_hd__and4_2 _26511_ (.A(iX[35]),
    .B(iX[36]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_16561_));
 sky130_fd_sc_hd__a22oi_2 _26512_ (.A1(iX[36]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[35]),
    .Y(_16562_));
 sky130_fd_sc_hd__nand2_2 _26513_ (.A(iX[34]),
    .B(iY[49]),
    .Y(_16564_));
 sky130_fd_sc_hd__o21a_2 _26514_ (.A1(_16561_),
    .A2(_16562_),
    .B1(_16564_),
    .X(_16565_));
 sky130_fd_sc_hd__nor3_2 _26515_ (.A(_16561_),
    .B(_16562_),
    .C(_16564_),
    .Y(_16566_));
 sky130_fd_sc_hd__nor2_2 _26516_ (.A(_16565_),
    .B(_16566_),
    .Y(_16567_));
 sky130_fd_sc_hd__xnor2_2 _26517_ (.A(_16560_),
    .B(_16567_),
    .Y(_16568_));
 sky130_fd_sc_hd__xnor2_2 _26518_ (.A(_16559_),
    .B(_16568_),
    .Y(_16569_));
 sky130_fd_sc_hd__a21o_2 _26519_ (.A1(_16558_),
    .A2(_16431_),
    .B1(_16569_),
    .X(_16570_));
 sky130_fd_sc_hd__nand3_2 _26520_ (.A(_16558_),
    .B(_16431_),
    .C(_16569_),
    .Y(_16571_));
 sky130_fd_sc_hd__nand2_2 _26521_ (.A(_16570_),
    .B(_16571_),
    .Y(_16572_));
 sky130_fd_sc_hd__or3_2 _26522_ (.A(_16556_),
    .B(_16557_),
    .C(_16572_),
    .X(_16573_));
 sky130_fd_sc_hd__o21ai_2 _26523_ (.A1(_16556_),
    .A2(_16557_),
    .B1(_16572_),
    .Y(_16575_));
 sky130_fd_sc_hd__and3_2 _26524_ (.A(_16555_),
    .B(_16573_),
    .C(_16575_),
    .X(_16576_));
 sky130_fd_sc_hd__a21oi_2 _26525_ (.A1(_16573_),
    .A2(_16575_),
    .B1(_16555_),
    .Y(_16577_));
 sky130_fd_sc_hd__nor2_2 _26526_ (.A(_16576_),
    .B(_16577_),
    .Y(_16578_));
 sky130_fd_sc_hd__o21a_2 _26527_ (.A1(_16554_),
    .A2(_16438_),
    .B1(_16578_),
    .X(_16579_));
 sky130_fd_sc_hd__or3_2 _26528_ (.A(_16554_),
    .B(_16438_),
    .C(_16578_),
    .X(_16580_));
 sky130_fd_sc_hd__or2b_2 _26529_ (.A(_16579_),
    .B_N(_16580_),
    .X(_16581_));
 sky130_fd_sc_hd__xnor2_2 _26530_ (.A(_16553_),
    .B(_16581_),
    .Y(_16582_));
 sky130_fd_sc_hd__or2b_2 _26531_ (.A(_16418_),
    .B_N(_16446_),
    .X(_16583_));
 sky130_fd_sc_hd__xnor2_2 _26532_ (.A(_16582_),
    .B(_16583_),
    .Y(_16584_));
 sky130_fd_sc_hd__a21o_2 _26533_ (.A1(_16420_),
    .A2(_16442_),
    .B1(_16440_),
    .X(_16586_));
 sky130_fd_sc_hd__xnor2_2 _26534_ (.A(_16584_),
    .B(_16586_),
    .Y(_16587_));
 sky130_fd_sc_hd__o21bai_2 _26535_ (.A1(_16447_),
    .A2(_16485_),
    .B1_N(_16587_),
    .Y(_16588_));
 sky130_fd_sc_hd__or3b_2 _26536_ (.A(_16447_),
    .B(_16485_),
    .C_N(_16587_),
    .X(_16589_));
 sky130_fd_sc_hd__nand3_2 _26537_ (.A(_16452_),
    .B(_16588_),
    .C(_16589_),
    .Y(_16590_));
 sky130_fd_sc_hd__a21o_2 _26538_ (.A1(_16588_),
    .A2(_16589_),
    .B1(_16452_),
    .X(_16591_));
 sky130_fd_sc_hd__and3_2 _26539_ (.A(_16455_),
    .B(_16590_),
    .C(_16591_),
    .X(_16592_));
 sky130_fd_sc_hd__a21oi_2 _26540_ (.A1(_16590_),
    .A2(_16591_),
    .B1(_16455_),
    .Y(_16593_));
 sky130_fd_sc_hd__or2_2 _26541_ (.A(_16592_),
    .B(_16593_),
    .X(_16594_));
 sky130_fd_sc_hd__or2b_2 _26542_ (.A(_16457_),
    .B_N(_16461_),
    .X(_16595_));
 sky130_fd_sc_hd__xnor2_2 _26543_ (.A(_16594_),
    .B(_16595_),
    .Y(_16597_));
 sky130_fd_sc_hd__nand2_2 _26544_ (.A(_16228_),
    .B(_16349_),
    .Y(_16598_));
 sky130_fd_sc_hd__nor2_2 _26545_ (.A(_16346_),
    .B(_16348_),
    .Y(_16599_));
 sky130_fd_sc_hd__and2b_2 _26546_ (.A_N(_16232_),
    .B(_16260_),
    .X(_16600_));
 sky130_fd_sc_hd__a31o_2 _26547_ (.A1(_15846_),
    .A2(_15845_),
    .A3(_16261_),
    .B1(_16600_),
    .X(_16601_));
 sky130_fd_sc_hd__nor2_2 _26548_ (.A(_16246_),
    .B(_16247_),
    .Y(_16602_));
 sky130_fd_sc_hd__a21o_2 _26549_ (.A1(_16248_),
    .A2(_16259_),
    .B1(_16602_),
    .X(_16603_));
 sky130_fd_sc_hd__and2b_2 _26550_ (.A_N(_16266_),
    .B(_16285_),
    .X(_16604_));
 sky130_fd_sc_hd__a21o_2 _26551_ (.A1(_16264_),
    .A2(_16286_),
    .B1(_16604_),
    .X(_16605_));
 sky130_fd_sc_hd__buf_1 _26552_ (.A(_16258_),
    .X(_16606_));
 sky130_fd_sc_hd__nand2_2 _26553_ (.A(iY[19]),
    .B(iY[51]),
    .Y(_16608_));
 sky130_fd_sc_hd__or2_2 _26554_ (.A(iY[19]),
    .B(iY[51]),
    .X(_16609_));
 sky130_fd_sc_hd__nand2_2 _26555_ (.A(_16608_),
    .B(_16609_),
    .Y(_16610_));
 sky130_fd_sc_hd__a21oi_2 _26556_ (.A1(_16251_),
    .A2(_16254_),
    .B1(_16249_),
    .Y(_16611_));
 sky130_fd_sc_hd__xor2_2 _26557_ (.A(_16610_),
    .B(_16611_),
    .X(_16612_));
 sky130_fd_sc_hd__buf_1 _26558_ (.A(_16612_),
    .X(_16613_));
 sky130_fd_sc_hd__buf_1 _26559_ (.A(_16613_),
    .X(_16614_));
 sky130_fd_sc_hd__a2bb2o_2 _26560_ (.A1_N(_11571_),
    .A2_N(_16606_),
    .B1(_16614_),
    .B2(_14592_),
    .X(_16615_));
 sky130_fd_sc_hd__xnor2_2 _26561_ (.A(_16610_),
    .B(_16611_),
    .Y(_16616_));
 sky130_fd_sc_hd__buf_1 _26562_ (.A(_16616_),
    .X(_16617_));
 sky130_fd_sc_hd__buf_1 _26563_ (.A(_16617_),
    .X(_16619_));
 sky130_fd_sc_hd__or3b_2 _26564_ (.A(_11571_),
    .B(_16619_),
    .C_N(_16259_),
    .X(_16620_));
 sky130_fd_sc_hd__nand2_2 _26565_ (.A(_16615_),
    .B(_16620_),
    .Y(_16621_));
 sky130_fd_sc_hd__nand2_2 _26566_ (.A(_16238_),
    .B(_16240_),
    .Y(_16622_));
 sky130_fd_sc_hd__or2_2 _26567_ (.A(_15858_),
    .B(_16269_),
    .X(_16623_));
 sky130_fd_sc_hd__a21bo_2 _26568_ (.A1(_16270_),
    .A2(_16272_),
    .B1_N(_16623_),
    .X(_16624_));
 sky130_fd_sc_hd__buf_1 _26569_ (.A(_12468_),
    .X(_16625_));
 sky130_fd_sc_hd__nor2_2 _26570_ (.A(_16625_),
    .B(_15835_),
    .Y(_16626_));
 sky130_fd_sc_hd__or4_2 _26571_ (.A(_15167_),
    .B(_14346_),
    .C(_16237_),
    .D(_15598_),
    .X(_16627_));
 sky130_fd_sc_hd__a2bb2o_2 _26572_ (.A1_N(_15167_),
    .A2_N(_15598_),
    .B1(_15585_),
    .B2(_14628_),
    .X(_16628_));
 sky130_fd_sc_hd__nand2_2 _26573_ (.A(_16627_),
    .B(_16628_),
    .Y(_16630_));
 sky130_fd_sc_hd__xnor2_2 _26574_ (.A(_16626_),
    .B(_16630_),
    .Y(_16631_));
 sky130_fd_sc_hd__xor2_2 _26575_ (.A(_16624_),
    .B(_16631_),
    .X(_16632_));
 sky130_fd_sc_hd__xor2_2 _26576_ (.A(_16622_),
    .B(_16632_),
    .X(_16633_));
 sky130_fd_sc_hd__a21o_2 _26577_ (.A1(_16233_),
    .A2(_16244_),
    .B1(_16242_),
    .X(_16634_));
 sky130_fd_sc_hd__xnor2_2 _26578_ (.A(_16633_),
    .B(_16634_),
    .Y(_16635_));
 sky130_fd_sc_hd__xnor2_2 _26579_ (.A(_16621_),
    .B(_16635_),
    .Y(_16636_));
 sky130_fd_sc_hd__xnor2_2 _26580_ (.A(_16605_),
    .B(_16636_),
    .Y(_16637_));
 sky130_fd_sc_hd__xnor2_2 _26581_ (.A(_16603_),
    .B(_16637_),
    .Y(_16638_));
 sky130_fd_sc_hd__o21ba_2 _26582_ (.A1(_16273_),
    .A2(_16284_),
    .B1_N(_16282_),
    .X(_16639_));
 sky130_fd_sc_hd__and2_2 _26583_ (.A(_16294_),
    .B(_16299_),
    .X(_16641_));
 sky130_fd_sc_hd__nand2_2 _26584_ (.A(_16277_),
    .B(_14608_),
    .Y(_16642_));
 sky130_fd_sc_hd__a22o_2 _26585_ (.A1(_16277_),
    .A2(_14410_),
    .B1(_14605_),
    .B2(_12816_),
    .X(_16643_));
 sky130_fd_sc_hd__o21a_2 _26586_ (.A1(_16269_),
    .A2(_16642_),
    .B1(_16643_),
    .X(_16644_));
 sky130_fd_sc_hd__nor2_2 _26587_ (.A(_14640_),
    .B(_14948_),
    .Y(_16645_));
 sky130_fd_sc_hd__xnor2_2 _26588_ (.A(_16644_),
    .B(_16645_),
    .Y(_16646_));
 sky130_fd_sc_hd__nand2_2 _26589_ (.A(_13845_),
    .B(_13887_),
    .Y(_16647_));
 sky130_fd_sc_hd__o22a_2 _26590_ (.A1(_14612_),
    .A2(_13842_),
    .B1(_13893_),
    .B2(_13502_),
    .X(_16648_));
 sky130_fd_sc_hd__o21ba_2 _26591_ (.A1(_16275_),
    .A2(_16647_),
    .B1_N(_16648_),
    .X(_16649_));
 sky130_fd_sc_hd__nand2_2 _26592_ (.A(_14652_),
    .B(_14392_),
    .Y(_16650_));
 sky130_fd_sc_hd__xor2_2 _26593_ (.A(_16649_),
    .B(_16650_),
    .X(_16652_));
 sky130_fd_sc_hd__o22a_2 _26594_ (.A1(_16274_),
    .A2(_16275_),
    .B1(_16276_),
    .B2(_16279_),
    .X(_16653_));
 sky130_fd_sc_hd__xnor2_2 _26595_ (.A(_16652_),
    .B(_16653_),
    .Y(_16654_));
 sky130_fd_sc_hd__xor2_2 _26596_ (.A(_16646_),
    .B(_16654_),
    .X(_16655_));
 sky130_fd_sc_hd__o21ai_2 _26597_ (.A1(_16641_),
    .A2(_16302_),
    .B1(_16655_),
    .Y(_16656_));
 sky130_fd_sc_hd__or3_2 _26598_ (.A(_16641_),
    .B(_16302_),
    .C(_16655_),
    .X(_16657_));
 sky130_fd_sc_hd__nand2_2 _26599_ (.A(_16656_),
    .B(_16657_),
    .Y(_16658_));
 sky130_fd_sc_hd__xor2_2 _26600_ (.A(_16639_),
    .B(_16658_),
    .X(_16659_));
 sky130_fd_sc_hd__a21bo_2 _26601_ (.A1(_16296_),
    .A2(_16298_),
    .B1_N(_16295_),
    .X(_16660_));
 sky130_fd_sc_hd__a21bo_2 _26602_ (.A1(_16305_),
    .A2(_16307_),
    .B1_N(_16306_),
    .X(_16661_));
 sky130_fd_sc_hd__nor2_2 _26603_ (.A(_12773_),
    .B(_14987_),
    .Y(_16663_));
 sky130_fd_sc_hd__o22a_2 _26604_ (.A1(_12850_),
    .A2(_14987_),
    .B1(_15004_),
    .B2(_12773_),
    .X(_16664_));
 sky130_fd_sc_hd__a31o_2 _26605_ (.A1(_14637_),
    .A2(_16292_),
    .A3(_16663_),
    .B1(_16664_),
    .X(_16665_));
 sky130_fd_sc_hd__nor2_2 _26606_ (.A(_14641_),
    .B(_15647_),
    .Y(_16666_));
 sky130_fd_sc_hd__xnor2_2 _26607_ (.A(_16665_),
    .B(_16666_),
    .Y(_16667_));
 sky130_fd_sc_hd__xor2_2 _26608_ (.A(_16661_),
    .B(_16667_),
    .X(_16668_));
 sky130_fd_sc_hd__xnor2_2 _26609_ (.A(_16660_),
    .B(_16668_),
    .Y(_16669_));
 sky130_fd_sc_hd__nor2_2 _26610_ (.A(_14356_),
    .B(_14998_),
    .Y(_16670_));
 sky130_fd_sc_hd__nor2_2 _26611_ (.A(_13926_),
    .B(_15668_),
    .Y(_16671_));
 sky130_fd_sc_hd__or4b_2 _26612_ (.A(_12248_),
    .B(_15219_),
    .C(_15220_),
    .D_N(_16671_),
    .X(_16672_));
 sky130_fd_sc_hd__a31o_2 _26613_ (.A1(_12243_),
    .A2(_15224_),
    .A3(_15226_),
    .B1(_16671_),
    .X(_16674_));
 sky130_fd_sc_hd__nand3_2 _26614_ (.A(_16670_),
    .B(_16672_),
    .C(_16674_),
    .Y(_16675_));
 sky130_fd_sc_hd__a21o_2 _26615_ (.A1(_16672_),
    .A2(_16674_),
    .B1(_16670_),
    .X(_16676_));
 sky130_fd_sc_hd__xnor2_2 _26616_ (.A(_15897_),
    .B(_15898_),
    .Y(_16677_));
 sky130_fd_sc_hd__xnor2_2 _26617_ (.A(iX[19]),
    .B(iX[51]),
    .Y(_16678_));
 sky130_fd_sc_hd__a22oi_2 _26618_ (.A1(iX[18]),
    .A2(iX[50]),
    .B1(_16316_),
    .B2(_16318_),
    .Y(_16679_));
 sky130_fd_sc_hd__xor2_2 _26619_ (.A(_16678_),
    .B(_16679_),
    .X(_16680_));
 sky130_fd_sc_hd__and3_2 _26620_ (.A(_11583_),
    .B(_16321_),
    .C(_16680_),
    .X(_16681_));
 sky130_fd_sc_hd__and2_2 _26621_ (.A(_16319_),
    .B(_16320_),
    .X(_16682_));
 sky130_fd_sc_hd__a22o_2 _26622_ (.A1(_11583_),
    .A2(_16682_),
    .B1(_16680_),
    .B2(_11380_),
    .X(_16683_));
 sky130_fd_sc_hd__or4b_4 _26623_ (.A(_11791_),
    .B(_16677_),
    .C(_16681_),
    .D_N(_16683_),
    .X(_16685_));
 sky130_fd_sc_hd__xnor2_2 _26624_ (.A(_16678_),
    .B(_16679_),
    .Y(_16686_));
 sky130_fd_sc_hd__or3b_2 _26625_ (.A(_11575_),
    .B(_16686_),
    .C_N(_16321_),
    .X(_16687_));
 sky130_fd_sc_hd__a22o_2 _26626_ (.A1(_15675_),
    .A2(_15900_),
    .B1(_16687_),
    .B2(_16683_),
    .X(_16688_));
 sky130_fd_sc_hd__nand2_2 _26627_ (.A(_16319_),
    .B(_16320_),
    .Y(_16689_));
 sky130_fd_sc_hd__or3_2 _26628_ (.A(_11566_),
    .B(_16314_),
    .C(_16689_),
    .X(_16690_));
 sky130_fd_sc_hd__a21bo_2 _26629_ (.A1(_16313_),
    .A2(_16323_),
    .B1_N(_16690_),
    .X(_16691_));
 sky130_fd_sc_hd__nand3_2 _26630_ (.A(_16685_),
    .B(_16688_),
    .C(_16691_),
    .Y(_16692_));
 sky130_fd_sc_hd__a21o_2 _26631_ (.A1(_16685_),
    .A2(_16688_),
    .B1(_16691_),
    .X(_16693_));
 sky130_fd_sc_hd__nand4_2 _26632_ (.A(_16675_),
    .B(_16676_),
    .C(_16692_),
    .D(_16693_),
    .Y(_16694_));
 sky130_fd_sc_hd__a22o_2 _26633_ (.A1(_16675_),
    .A2(_16676_),
    .B1(_16692_),
    .B2(_16693_),
    .X(_16696_));
 sky130_fd_sc_hd__a31o_2 _26634_ (.A1(_16308_),
    .A2(_16309_),
    .A3(_16326_),
    .B1(_16325_),
    .X(_16697_));
 sky130_fd_sc_hd__and3_2 _26635_ (.A(_16694_),
    .B(_16696_),
    .C(_16697_),
    .X(_16698_));
 sky130_fd_sc_hd__a21oi_2 _26636_ (.A1(_16694_),
    .A2(_16696_),
    .B1(_16697_),
    .Y(_16699_));
 sky130_fd_sc_hd__nor3_2 _26637_ (.A(_16669_),
    .B(_16698_),
    .C(_16699_),
    .Y(_16700_));
 sky130_fd_sc_hd__o21a_2 _26638_ (.A1(_16698_),
    .A2(_16699_),
    .B1(_16669_),
    .X(_16701_));
 sky130_fd_sc_hd__or2_2 _26639_ (.A(_16700_),
    .B(_16701_),
    .X(_16702_));
 sky130_fd_sc_hd__o32a_2 _26640_ (.A1(_16302_),
    .A2(_16303_),
    .A3(_16331_),
    .B1(_16330_),
    .B2(_16328_),
    .X(_16703_));
 sky130_fd_sc_hd__xor2_2 _26641_ (.A(_16702_),
    .B(_16703_),
    .X(_16704_));
 sky130_fd_sc_hd__xor2_2 _26642_ (.A(_16659_),
    .B(_16704_),
    .X(_16705_));
 sky130_fd_sc_hd__nand2_2 _26643_ (.A(_16332_),
    .B(_16335_),
    .Y(_16707_));
 sky130_fd_sc_hd__a21bo_2 _26644_ (.A1(_16287_),
    .A2(_16336_),
    .B1_N(_16707_),
    .X(_16708_));
 sky130_fd_sc_hd__xnor2_2 _26645_ (.A(_16705_),
    .B(_16708_),
    .Y(_16709_));
 sky130_fd_sc_hd__xnor2_2 _26646_ (.A(_16638_),
    .B(_16709_),
    .Y(_16710_));
 sky130_fd_sc_hd__or2b_2 _26647_ (.A(_16339_),
    .B_N(_16337_),
    .X(_16711_));
 sky130_fd_sc_hd__a21bo_2 _26648_ (.A1(_16262_),
    .A2(_16340_),
    .B1_N(_16711_),
    .X(_16712_));
 sky130_fd_sc_hd__xnor2_2 _26649_ (.A(_16710_),
    .B(_16712_),
    .Y(_16713_));
 sky130_fd_sc_hd__xnor2_2 _26650_ (.A(_16601_),
    .B(_16713_),
    .Y(_16714_));
 sky130_fd_sc_hd__nor2_2 _26651_ (.A(_16341_),
    .B(_16343_),
    .Y(_16715_));
 sky130_fd_sc_hd__a21oi_2 _26652_ (.A1(_16229_),
    .A2(_16345_),
    .B1(_16715_),
    .Y(_16716_));
 sky130_fd_sc_hd__xor2_2 _26653_ (.A(_16714_),
    .B(_16716_),
    .X(_16718_));
 sky130_fd_sc_hd__xnor2_2 _26654_ (.A(_16599_),
    .B(_16718_),
    .Y(_16719_));
 sky130_fd_sc_hd__xor2_2 _26655_ (.A(_16598_),
    .B(_16719_),
    .X(_16720_));
 sky130_fd_sc_hd__a32o_2 _26656_ (.A1(_15823_),
    .A2(_15926_),
    .A3(_16350_),
    .B1(_16351_),
    .B2(_16353_),
    .X(_16721_));
 sky130_fd_sc_hd__xnor2_2 _26657_ (.A(_16720_),
    .B(_16721_),
    .Y(_16722_));
 sky130_fd_sc_hd__xnor2_2 _26658_ (.A(_16597_),
    .B(_16722_),
    .Y(_16723_));
 sky130_fd_sc_hd__xnor2_2 _26659_ (.A(oO[19]),
    .B(_16723_),
    .Y(_16724_));
 sky130_fd_sc_hd__or2b_2 _26660_ (.A(_16354_),
    .B_N(_16463_),
    .X(_16725_));
 sky130_fd_sc_hd__o21a_2 _26661_ (.A1(oO[18]),
    .A2(_16464_),
    .B1(_16725_),
    .X(_16726_));
 sky130_fd_sc_hd__xor2_2 _26662_ (.A(_16724_),
    .B(_16726_),
    .X(_16727_));
 sky130_fd_sc_hd__nand2_2 _26663_ (.A(_16475_),
    .B(_16727_),
    .Y(_16729_));
 sky130_fd_sc_hd__or3b_2 _26664_ (.A(_16469_),
    .B(_16727_),
    .C_N(_16466_),
    .X(_16730_));
 sky130_fd_sc_hd__a311o_2 _26665_ (.A1(_16471_),
    .A2(_16472_),
    .A3(_16473_),
    .B1(_16727_),
    .C1(_16470_),
    .X(_16731_));
 sky130_fd_sc_hd__and2_2 _26666_ (.A(_16730_),
    .B(_16731_),
    .X(_16732_));
 sky130_fd_sc_hd__o21ai_2 _26667_ (.A1(_16484_),
    .A2(_16729_),
    .B1(_16732_),
    .Y(_16733_));
 sky130_fd_sc_hd__and2b_2 _26668_ (.A_N(_16216_),
    .B(_16215_),
    .X(_16734_));
 sky130_fd_sc_hd__and3b_2 _26669_ (.A_N(_15487_),
    .B(iX[31]),
    .C(iY[20]),
    .X(_16735_));
 sky130_fd_sc_hd__and2_2 _26670_ (.A(iY[22]),
    .B(iX[30]),
    .X(_16736_));
 sky130_fd_sc_hd__and3_2 _26671_ (.A(iY[21]),
    .B(iX[29]),
    .C(_16736_),
    .X(_16737_));
 sky130_fd_sc_hd__a22oi_2 _26672_ (.A1(iY[22]),
    .A2(iX[29]),
    .B1(iX[30]),
    .B2(iY[21]),
    .Y(_16738_));
 sky130_fd_sc_hd__and4bb_2 _26673_ (.A_N(_16737_),
    .B_N(_16738_),
    .C(iY[23]),
    .D(iX[28]),
    .X(_16740_));
 sky130_fd_sc_hd__o2bb2a_2 _26674_ (.A1_N(iY[23]),
    .A2_N(iX[28]),
    .B1(_16737_),
    .B2(_16738_),
    .X(_16741_));
 sky130_fd_sc_hd__nor2_2 _26675_ (.A(_16740_),
    .B(_16741_),
    .Y(_16742_));
 sky130_fd_sc_hd__xnor2_2 _26676_ (.A(_16735_),
    .B(_16742_),
    .Y(_16743_));
 sky130_fd_sc_hd__or2b_2 _26677_ (.A(_16167_),
    .B_N(_16166_),
    .X(_16744_));
 sky130_fd_sc_hd__and4_2 _26678_ (.A(iX[23]),
    .B(iX[24]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_16745_));
 sky130_fd_sc_hd__a22oi_2 _26679_ (.A1(iX[24]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[23]),
    .Y(_16746_));
 sky130_fd_sc_hd__nor2_2 _26680_ (.A(_16745_),
    .B(_16746_),
    .Y(_16747_));
 sky130_fd_sc_hd__nand2_2 _26681_ (.A(iX[22]),
    .B(iY[29]),
    .Y(_16748_));
 sky130_fd_sc_hd__xnor2_2 _26682_ (.A(_16747_),
    .B(_16748_),
    .Y(_16749_));
 sky130_fd_sc_hd__o21ba_2 _26683_ (.A1(_16163_),
    .A2(_16165_),
    .B1_N(_16162_),
    .X(_16751_));
 sky130_fd_sc_hd__xnor2_2 _26684_ (.A(_16749_),
    .B(_16751_),
    .Y(_16752_));
 sky130_fd_sc_hd__nand3_2 _26685_ (.A(iX[21]),
    .B(iY[30]),
    .C(_16752_),
    .Y(_16753_));
 sky130_fd_sc_hd__a21o_2 _26686_ (.A1(iX[21]),
    .A2(iY[30]),
    .B1(_16752_),
    .X(_16754_));
 sky130_fd_sc_hd__nand2_2 _26687_ (.A(_16753_),
    .B(_16754_),
    .Y(_16755_));
 sky130_fd_sc_hd__a21oi_2 _26688_ (.A1(_16744_),
    .A2(_16172_),
    .B1(_16755_),
    .Y(_16756_));
 sky130_fd_sc_hd__and3_2 _26689_ (.A(_16744_),
    .B(_16172_),
    .C(_16755_),
    .X(_16757_));
 sky130_fd_sc_hd__nor2_2 _26690_ (.A(_16756_),
    .B(_16757_),
    .Y(_16758_));
 sky130_fd_sc_hd__nand2_2 _26691_ (.A(iX[20]),
    .B(iY[31]),
    .Y(_16759_));
 sky130_fd_sc_hd__xnor2_2 _26692_ (.A(_16758_),
    .B(_16759_),
    .Y(_16760_));
 sky130_fd_sc_hd__or2b_2 _26693_ (.A(_16183_),
    .B_N(_16192_),
    .X(_16762_));
 sky130_fd_sc_hd__or2b_2 _26694_ (.A(_16144_),
    .B_N(_16145_),
    .X(_16763_));
 sky130_fd_sc_hd__o21ba_2 _26695_ (.A1(_16149_),
    .A2(_16151_),
    .B1_N(_16148_),
    .X(_16764_));
 sky130_fd_sc_hd__and4_2 _26696_ (.A(iY[24]),
    .B(iY[25]),
    .C(iX[26]),
    .D(iX[27]),
    .X(_16765_));
 sky130_fd_sc_hd__a22oi_2 _26697_ (.A1(iY[25]),
    .A2(iX[26]),
    .B1(iX[27]),
    .B2(iY[24]),
    .Y(_16766_));
 sky130_fd_sc_hd__nor2_2 _26698_ (.A(_16765_),
    .B(_16766_),
    .Y(_16767_));
 sky130_fd_sc_hd__nand2_2 _26699_ (.A(iX[25]),
    .B(iY[26]),
    .Y(_16768_));
 sky130_fd_sc_hd__xnor2_2 _26700_ (.A(_16767_),
    .B(_16768_),
    .Y(_16769_));
 sky130_fd_sc_hd__xnor2_2 _26701_ (.A(_16764_),
    .B(_16769_),
    .Y(_16770_));
 sky130_fd_sc_hd__o21a_2 _26702_ (.A1(_16184_),
    .A2(_16186_),
    .B1(_16770_),
    .X(_16771_));
 sky130_fd_sc_hd__nor3_2 _26703_ (.A(_16184_),
    .B(_16186_),
    .C(_16770_),
    .Y(_16773_));
 sky130_fd_sc_hd__or2_2 _26704_ (.A(_16771_),
    .B(_16773_),
    .X(_16774_));
 sky130_fd_sc_hd__a21oi_2 _26705_ (.A1(_16763_),
    .A2(_16153_),
    .B1(_16774_),
    .Y(_16775_));
 sky130_fd_sc_hd__and3_2 _26706_ (.A(_16763_),
    .B(_16153_),
    .C(_16774_),
    .X(_16776_));
 sky130_fd_sc_hd__a211o_2 _26707_ (.A1(_16189_),
    .A2(_16762_),
    .B1(_16775_),
    .C1(_16776_),
    .X(_16777_));
 sky130_fd_sc_hd__o211ai_2 _26708_ (.A1(_16775_),
    .A2(_16776_),
    .B1(_16189_),
    .C1(_16762_),
    .Y(_16778_));
 sky130_fd_sc_hd__o211ai_2 _26709_ (.A1(_16194_),
    .A2(_16196_),
    .B1(_16777_),
    .C1(_16778_),
    .Y(_16779_));
 sky130_fd_sc_hd__a211o_2 _26710_ (.A1(_16777_),
    .A2(_16778_),
    .B1(_16194_),
    .C1(_16196_),
    .X(_16780_));
 sky130_fd_sc_hd__and3_2 _26711_ (.A(_16760_),
    .B(_16779_),
    .C(_16780_),
    .X(_16781_));
 sky130_fd_sc_hd__a21oi_2 _26712_ (.A1(_16779_),
    .A2(_16780_),
    .B1(_16760_),
    .Y(_16782_));
 sky130_fd_sc_hd__nor3_2 _26713_ (.A(_16156_),
    .B(_16781_),
    .C(_16782_),
    .Y(_16784_));
 sky130_fd_sc_hd__o21a_2 _26714_ (.A1(_16781_),
    .A2(_16782_),
    .B1(_16156_),
    .X(_16785_));
 sky130_fd_sc_hd__a211oi_2 _26715_ (.A1(_16199_),
    .A2(_16202_),
    .B1(_16784_),
    .C1(_16785_),
    .Y(_16786_));
 sky130_fd_sc_hd__o211a_2 _26716_ (.A1(_16784_),
    .A2(_16785_),
    .B1(_16199_),
    .C1(_16202_),
    .X(_16787_));
 sky130_fd_sc_hd__or3_2 _26717_ (.A(_16743_),
    .B(_16786_),
    .C(_16787_),
    .X(_16788_));
 sky130_fd_sc_hd__o21ai_2 _26718_ (.A1(_16786_),
    .A2(_16787_),
    .B1(_16743_),
    .Y(_16789_));
 sky130_fd_sc_hd__and3_2 _26719_ (.A(_16208_),
    .B(_16788_),
    .C(_16789_),
    .X(_16790_));
 sky130_fd_sc_hd__a21oi_2 _26720_ (.A1(_16788_),
    .A2(_16789_),
    .B1(_16208_),
    .Y(_16791_));
 sky130_fd_sc_hd__nor2_2 _26721_ (.A(_16790_),
    .B(_16791_),
    .Y(_16792_));
 sky130_fd_sc_hd__o21a_2 _26722_ (.A1(_16204_),
    .A2(_16206_),
    .B1(_16792_),
    .X(_16793_));
 sky130_fd_sc_hd__nor3_2 _26723_ (.A(_16204_),
    .B(_16206_),
    .C(_16792_),
    .Y(_16795_));
 sky130_fd_sc_hd__a211oi_2 _26724_ (.A1(_16210_),
    .A2(_16213_),
    .B1(_16793_),
    .C1(_16795_),
    .Y(_16796_));
 sky130_fd_sc_hd__o211a_2 _26725_ (.A1(_16793_),
    .A2(_16795_),
    .B1(_16210_),
    .C1(_16213_),
    .X(_16797_));
 sky130_fd_sc_hd__nor2_2 _26726_ (.A(_16796_),
    .B(_16797_),
    .Y(_16798_));
 sky130_fd_sc_hd__a31o_2 _26727_ (.A1(iX[19]),
    .A2(iY[31]),
    .A3(_16176_),
    .B1(_16174_),
    .X(_16799_));
 sky130_fd_sc_hd__xor2_2 _26728_ (.A(_16798_),
    .B(_16799_),
    .X(_16800_));
 sky130_fd_sc_hd__or3_2 _26729_ (.A(_16734_),
    .B(_16218_),
    .C(_16800_),
    .X(_16801_));
 sky130_fd_sc_hd__inv_2 _26730_ (.A(_16801_),
    .Y(_16802_));
 sky130_fd_sc_hd__o21a_2 _26731_ (.A1(_16734_),
    .A2(_16218_),
    .B1(_16800_),
    .X(_16803_));
 sky130_fd_sc_hd__nor2_2 _26732_ (.A(_16802_),
    .B(_16803_),
    .Y(_16804_));
 sky130_fd_sc_hd__and2b_2 _26733_ (.A_N(_16221_),
    .B(_16220_),
    .X(_16806_));
 sky130_fd_sc_hd__and2b_2 _26734_ (.A_N(_16225_),
    .B(_16222_),
    .X(_16807_));
 sky130_fd_sc_hd__nor2_2 _26735_ (.A(_16806_),
    .B(_16807_),
    .Y(_16808_));
 sky130_fd_sc_hd__xor2_2 _26736_ (.A(_16804_),
    .B(_16808_),
    .X(_16809_));
 sky130_fd_sc_hd__and2_2 _26737_ (.A(_16733_),
    .B(_16809_),
    .X(_16810_));
 sky130_fd_sc_hd__nor2_2 _26738_ (.A(_16733_),
    .B(_16809_),
    .Y(_16811_));
 sky130_fd_sc_hd__nor2_2 _26739_ (.A(_16810_),
    .B(_16811_),
    .Y(_16812_));
 sky130_fd_sc_hd__a21oi_2 _26740_ (.A1(_16480_),
    .A2(_16483_),
    .B1(_16478_),
    .Y(_16813_));
 sky130_fd_sc_hd__xnor2_2 _26741_ (.A(_16812_),
    .B(_16813_),
    .Y(oO[51]));
 sky130_fd_sc_hd__and2_2 _26742_ (.A(_16222_),
    .B(_16804_),
    .X(_16814_));
 sky130_fd_sc_hd__and2b_2 _26743_ (.A_N(_16224_),
    .B(_16814_),
    .X(_16816_));
 sky130_fd_sc_hd__o2111a_2 _26744_ (.A1(_15473_),
    .A2(_15476_),
    .B1(_15572_),
    .C1(_16132_),
    .D1(_16814_),
    .X(_16817_));
 sky130_fd_sc_hd__a21o_2 _26745_ (.A1(_16806_),
    .A2(_16801_),
    .B1(_16803_),
    .X(_16818_));
 sky130_fd_sc_hd__and3_2 _26746_ (.A(iY[21]),
    .B(iX[31]),
    .C(_16736_),
    .X(_16819_));
 sky130_fd_sc_hd__a21o_2 _26747_ (.A1(iY[21]),
    .A2(iX[31]),
    .B1(_16736_),
    .X(_16820_));
 sky130_fd_sc_hd__and2b_2 _26748_ (.A_N(_16819_),
    .B(_16820_),
    .X(_16821_));
 sky130_fd_sc_hd__nand2_2 _26749_ (.A(iY[23]),
    .B(iX[29]),
    .Y(_16822_));
 sky130_fd_sc_hd__xnor2_2 _26750_ (.A(_16821_),
    .B(_16822_),
    .Y(_16823_));
 sky130_fd_sc_hd__inv_2 _26751_ (.A(_16823_),
    .Y(_16824_));
 sky130_fd_sc_hd__inv_2 _26752_ (.A(_16781_),
    .Y(_16825_));
 sky130_fd_sc_hd__a21o_2 _26753_ (.A1(_16763_),
    .A2(_16153_),
    .B1(_16774_),
    .X(_16827_));
 sky130_fd_sc_hd__and2b_2 _26754_ (.A_N(_16764_),
    .B(_16769_),
    .X(_16828_));
 sky130_fd_sc_hd__a21oi_2 _26755_ (.A1(_16735_),
    .A2(_16742_),
    .B1(_16142_),
    .Y(_16829_));
 sky130_fd_sc_hd__o21ba_2 _26756_ (.A1(_16766_),
    .A2(_16768_),
    .B1_N(_16765_),
    .X(_16830_));
 sky130_fd_sc_hd__and4_2 _26757_ (.A(iY[24]),
    .B(iY[25]),
    .C(iX[27]),
    .D(iX[28]),
    .X(_16831_));
 sky130_fd_sc_hd__a22oi_2 _26758_ (.A1(iY[25]),
    .A2(iX[27]),
    .B1(iX[28]),
    .B2(iY[24]),
    .Y(_16832_));
 sky130_fd_sc_hd__nor2_2 _26759_ (.A(_16831_),
    .B(_16832_),
    .Y(_16833_));
 sky130_fd_sc_hd__nand2_2 _26760_ (.A(iX[26]),
    .B(iY[26]),
    .Y(_16834_));
 sky130_fd_sc_hd__xnor2_2 _26761_ (.A(_16833_),
    .B(_16834_),
    .Y(_16835_));
 sky130_fd_sc_hd__o21a_2 _26762_ (.A1(_16737_),
    .A2(_16740_),
    .B1(_16835_),
    .X(_16836_));
 sky130_fd_sc_hd__nor3_2 _26763_ (.A(_16737_),
    .B(_16740_),
    .C(_16835_),
    .Y(_16838_));
 sky130_fd_sc_hd__nor2_2 _26764_ (.A(_16836_),
    .B(_16838_),
    .Y(_16839_));
 sky130_fd_sc_hd__xnor2_2 _26765_ (.A(_16830_),
    .B(_16839_),
    .Y(_16840_));
 sky130_fd_sc_hd__xnor2_2 _26766_ (.A(_16829_),
    .B(_16840_),
    .Y(_16841_));
 sky130_fd_sc_hd__o21a_2 _26767_ (.A1(_16828_),
    .A2(_16771_),
    .B1(_16841_),
    .X(_16842_));
 sky130_fd_sc_hd__nor3_2 _26768_ (.A(_16828_),
    .B(_16771_),
    .C(_16841_),
    .Y(_16843_));
 sky130_fd_sc_hd__a211oi_2 _26769_ (.A1(_16827_),
    .A2(_16777_),
    .B1(_16842_),
    .C1(_16843_),
    .Y(_16844_));
 sky130_fd_sc_hd__inv_2 _26770_ (.A(_16844_),
    .Y(_16845_));
 sky130_fd_sc_hd__o211ai_2 _26771_ (.A1(_16842_),
    .A2(_16843_),
    .B1(_16827_),
    .C1(_16777_),
    .Y(_16846_));
 sky130_fd_sc_hd__or2b_2 _26772_ (.A(_16751_),
    .B_N(_16749_),
    .X(_16847_));
 sky130_fd_sc_hd__and4_2 _26773_ (.A(iX[24]),
    .B(iX[25]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_16849_));
 sky130_fd_sc_hd__a22oi_2 _26774_ (.A1(iX[25]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[24]),
    .Y(_16850_));
 sky130_fd_sc_hd__nor2_2 _26775_ (.A(_16849_),
    .B(_16850_),
    .Y(_16851_));
 sky130_fd_sc_hd__nand2_2 _26776_ (.A(iX[23]),
    .B(iY[29]),
    .Y(_16852_));
 sky130_fd_sc_hd__xnor2_2 _26777_ (.A(_16851_),
    .B(_16852_),
    .Y(_16853_));
 sky130_fd_sc_hd__o21ba_2 _26778_ (.A1(_16746_),
    .A2(_16748_),
    .B1_N(_16745_),
    .X(_16854_));
 sky130_fd_sc_hd__xnor2_2 _26779_ (.A(_16853_),
    .B(_16854_),
    .Y(_16855_));
 sky130_fd_sc_hd__nand3_2 _26780_ (.A(iX[22]),
    .B(iY[30]),
    .C(_16855_),
    .Y(_16856_));
 sky130_fd_sc_hd__a21o_2 _26781_ (.A1(iX[22]),
    .A2(iY[30]),
    .B1(_16855_),
    .X(_16857_));
 sky130_fd_sc_hd__nand2_2 _26782_ (.A(_16856_),
    .B(_16857_),
    .Y(_16858_));
 sky130_fd_sc_hd__a21oi_2 _26783_ (.A1(_16847_),
    .A2(_16753_),
    .B1(_16858_),
    .Y(_16860_));
 sky130_fd_sc_hd__and3_2 _26784_ (.A(_16847_),
    .B(_16753_),
    .C(_16858_),
    .X(_16861_));
 sky130_fd_sc_hd__nor2_2 _26785_ (.A(_16860_),
    .B(_16861_),
    .Y(_16862_));
 sky130_fd_sc_hd__nand2_2 _26786_ (.A(iX[21]),
    .B(iY[31]),
    .Y(_16863_));
 sky130_fd_sc_hd__xnor2_2 _26787_ (.A(_16862_),
    .B(_16863_),
    .Y(_16864_));
 sky130_fd_sc_hd__and3_2 _26788_ (.A(_16845_),
    .B(_16846_),
    .C(_16864_),
    .X(_16865_));
 sky130_fd_sc_hd__a21oi_2 _26789_ (.A1(_16845_),
    .A2(_16846_),
    .B1(_16864_),
    .Y(_16866_));
 sky130_fd_sc_hd__a211o_2 _26790_ (.A1(_16779_),
    .A2(_16825_),
    .B1(_16865_),
    .C1(_16866_),
    .X(_16867_));
 sky130_fd_sc_hd__o211ai_2 _26791_ (.A1(_16865_),
    .A2(_16866_),
    .B1(_16779_),
    .C1(_16825_),
    .Y(_16868_));
 sky130_fd_sc_hd__nand2_2 _26792_ (.A(_16867_),
    .B(_16868_),
    .Y(_16869_));
 sky130_fd_sc_hd__nor2_2 _26793_ (.A(_16824_),
    .B(_16869_),
    .Y(_16871_));
 sky130_fd_sc_hd__and2_2 _26794_ (.A(_16824_),
    .B(_16869_),
    .X(_16872_));
 sky130_fd_sc_hd__or2_2 _26795_ (.A(_16871_),
    .B(_16872_),
    .X(_16873_));
 sky130_fd_sc_hd__or2_2 _26796_ (.A(_16788_),
    .B(_16873_),
    .X(_16874_));
 sky130_fd_sc_hd__nand2_2 _26797_ (.A(_16788_),
    .B(_16873_),
    .Y(_16875_));
 sky130_fd_sc_hd__and2_2 _26798_ (.A(_16874_),
    .B(_16875_),
    .X(_16876_));
 sky130_fd_sc_hd__o21ai_2 _26799_ (.A1(_16784_),
    .A2(_16786_),
    .B1(_16876_),
    .Y(_16877_));
 sky130_fd_sc_hd__or3_2 _26800_ (.A(_16784_),
    .B(_16786_),
    .C(_16876_),
    .X(_16878_));
 sky130_fd_sc_hd__and2_2 _26801_ (.A(_16877_),
    .B(_16878_),
    .X(_16879_));
 sky130_fd_sc_hd__o21ai_2 _26802_ (.A1(_16790_),
    .A2(_16793_),
    .B1(_16879_),
    .Y(_16880_));
 sky130_fd_sc_hd__or3_2 _26803_ (.A(_16790_),
    .B(_16793_),
    .C(_16879_),
    .X(_16882_));
 sky130_fd_sc_hd__nand2_2 _26804_ (.A(_16880_),
    .B(_16882_),
    .Y(_16883_));
 sky130_fd_sc_hd__a31o_2 _26805_ (.A1(iX[20]),
    .A2(iY[31]),
    .A3(_16758_),
    .B1(_16756_),
    .X(_16884_));
 sky130_fd_sc_hd__xnor2_2 _26806_ (.A(_16883_),
    .B(_16884_),
    .Y(_16885_));
 sky130_fd_sc_hd__a21oi_2 _26807_ (.A1(_16798_),
    .A2(_16799_),
    .B1(_16796_),
    .Y(_16886_));
 sky130_fd_sc_hd__xnor2_2 _26808_ (.A(_16885_),
    .B(_16886_),
    .Y(_16887_));
 sky130_fd_sc_hd__o31a_2 _26809_ (.A1(_16816_),
    .A2(_16817_),
    .A3(_16818_),
    .B1(_16887_),
    .X(_16888_));
 sky130_fd_sc_hd__or4_2 _26810_ (.A(_16816_),
    .B(_16817_),
    .C(_16818_),
    .D(_16887_),
    .X(_16889_));
 sky130_fd_sc_hd__nand2b_2 _26811_ (.A_N(_16888_),
    .B(_16889_),
    .Y(_16890_));
 sky130_fd_sc_hd__or2b_2 _26812_ (.A(_16726_),
    .B_N(_16724_),
    .X(_16891_));
 sky130_fd_sc_hd__and2_2 _26813_ (.A(_16351_),
    .B(_16720_),
    .X(_16893_));
 sky130_fd_sc_hd__and2_2 _26814_ (.A(_15710_),
    .B(_15927_),
    .X(_16894_));
 sky130_fd_sc_hd__nand2_2 _26815_ (.A(_16599_),
    .B(_16718_),
    .Y(_16895_));
 sky130_fd_sc_hd__or2_2 _26816_ (.A(_16599_),
    .B(_16718_),
    .X(_16896_));
 sky130_fd_sc_hd__and4b_2 _26817_ (.A_N(_16227_),
    .B(_16350_),
    .C(_16895_),
    .D(_16896_),
    .X(_16897_));
 sky130_fd_sc_hd__nor2_2 _26818_ (.A(_16598_),
    .B(_16719_),
    .Y(_16898_));
 sky130_fd_sc_hd__a311o_2 _26819_ (.A1(_16351_),
    .A2(_16352_),
    .A3(_16720_),
    .B1(_16897_),
    .C1(_16898_),
    .X(_16899_));
 sky130_fd_sc_hd__a31o_2 _26820_ (.A1(_15579_),
    .A2(_16893_),
    .A3(_16894_),
    .B1(_16899_),
    .X(_16900_));
 sky130_fd_sc_hd__nor2_2 _26821_ (.A(_16714_),
    .B(_16716_),
    .Y(_16901_));
 sky130_fd_sc_hd__or2b_2 _26822_ (.A(_16636_),
    .B_N(_16605_),
    .X(_16902_));
 sky130_fd_sc_hd__a21bo_2 _26823_ (.A1(_16603_),
    .A2(_16637_),
    .B1_N(_16902_),
    .X(_16904_));
 sky130_fd_sc_hd__o2bb2a_2 _26824_ (.A1_N(_16633_),
    .A2_N(_16634_),
    .B1(_16635_),
    .B2(_16621_),
    .X(_16905_));
 sky130_fd_sc_hd__o21ai_2 _26825_ (.A1(_16639_),
    .A2(_16658_),
    .B1(_16656_),
    .Y(_16906_));
 sky130_fd_sc_hd__nor2_2 _26826_ (.A(_12468_),
    .B(_16255_),
    .Y(_16907_));
 sky130_fd_sc_hd__or3b_2 _26827_ (.A(_11570_),
    .B(_16617_),
    .C_N(_16907_),
    .X(_16908_));
 sky130_fd_sc_hd__a21o_2 _26828_ (.A1(_12838_),
    .A2(_16613_),
    .B1(_16907_),
    .X(_16909_));
 sky130_fd_sc_hd__inv_2 _26829_ (.A(_15595_),
    .Y(_16910_));
 sky130_fd_sc_hd__or3_2 _26830_ (.A(_16249_),
    .B(_16250_),
    .C(_16610_),
    .X(_16911_));
 sky130_fd_sc_hd__or4b_4 _26831_ (.A(_16910_),
    .B(_15832_),
    .C(_16911_),
    .D_N(_15592_),
    .X(_16912_));
 sky130_fd_sc_hd__inv_2 _26832_ (.A(_16911_),
    .Y(_16913_));
 sky130_fd_sc_hd__a21bo_2 _26833_ (.A1(_16253_),
    .A2(_16913_),
    .B1_N(_16608_),
    .X(_16915_));
 sky130_fd_sc_hd__a21oi_2 _26834_ (.A1(_16249_),
    .A2(_16609_),
    .B1(_16915_),
    .Y(_16916_));
 sky130_fd_sc_hd__nand2_2 _26835_ (.A(_16912_),
    .B(_16916_),
    .Y(_16917_));
 sky130_fd_sc_hd__nand2_2 _26836_ (.A(iY[20]),
    .B(iY[52]),
    .Y(_16918_));
 sky130_fd_sc_hd__or2_2 _26837_ (.A(iY[20]),
    .B(iY[52]),
    .X(_16919_));
 sky130_fd_sc_hd__nand2_2 _26838_ (.A(_16918_),
    .B(_16919_),
    .Y(_16920_));
 sky130_fd_sc_hd__xor2_2 _26839_ (.A(_16917_),
    .B(_16920_),
    .X(_16921_));
 sky130_fd_sc_hd__buf_1 _26840_ (.A(_16921_),
    .X(_16922_));
 sky130_fd_sc_hd__nor2_2 _26841_ (.A(_11578_),
    .B(_16922_),
    .Y(_16923_));
 sky130_fd_sc_hd__and3_2 _26842_ (.A(_16908_),
    .B(_16909_),
    .C(_16923_),
    .X(_16924_));
 sky130_fd_sc_hd__a21oi_2 _26843_ (.A1(_16908_),
    .A2(_16909_),
    .B1(_16923_),
    .Y(_16926_));
 sky130_fd_sc_hd__or2_2 _26844_ (.A(_16924_),
    .B(_16926_),
    .X(_16927_));
 sky130_fd_sc_hd__nor2_2 _26845_ (.A(_16620_),
    .B(_16927_),
    .Y(_16928_));
 sky130_fd_sc_hd__and2_2 _26846_ (.A(_16620_),
    .B(_16927_),
    .X(_16929_));
 sky130_fd_sc_hd__nor2_2 _26847_ (.A(_16928_),
    .B(_16929_),
    .Y(_16930_));
 sky130_fd_sc_hd__a21bo_2 _26848_ (.A1(_16626_),
    .A2(_16628_),
    .B1_N(_16627_),
    .X(_16931_));
 sky130_fd_sc_hd__a2bb2o_2 _26849_ (.A1_N(_16269_),
    .A2_N(_16642_),
    .B1(_16643_),
    .B2(_16645_),
    .X(_16932_));
 sky130_fd_sc_hd__inv_2 _26850_ (.A(_15834_),
    .Y(_16933_));
 sky130_fd_sc_hd__buf_1 _26851_ (.A(_16933_),
    .X(_16934_));
 sky130_fd_sc_hd__or4_2 _26852_ (.A(_14346_),
    .B(_12457_),
    .C(_15153_),
    .D(_15597_),
    .X(_16935_));
 sky130_fd_sc_hd__a2bb2o_2 _26853_ (.A1_N(_14346_),
    .A2_N(_15597_),
    .B1(_15585_),
    .B2(_15624_),
    .X(_16937_));
 sky130_fd_sc_hd__nand4_2 _26854_ (.A(_14388_),
    .B(_16934_),
    .C(_16935_),
    .D(_16937_),
    .Y(_16938_));
 sky130_fd_sc_hd__a22o_2 _26855_ (.A1(_14388_),
    .A2(_16933_),
    .B1(_16935_),
    .B2(_16937_),
    .X(_16939_));
 sky130_fd_sc_hd__nand3_2 _26856_ (.A(_16932_),
    .B(_16938_),
    .C(_16939_),
    .Y(_16940_));
 sky130_fd_sc_hd__a21o_2 _26857_ (.A1(_16938_),
    .A2(_16939_),
    .B1(_16932_),
    .X(_16941_));
 sky130_fd_sc_hd__and3_2 _26858_ (.A(_16931_),
    .B(_16940_),
    .C(_16941_),
    .X(_16942_));
 sky130_fd_sc_hd__a21oi_2 _26859_ (.A1(_16940_),
    .A2(_16941_),
    .B1(_16931_),
    .Y(_16943_));
 sky130_fd_sc_hd__or2_2 _26860_ (.A(_16942_),
    .B(_16943_),
    .X(_16944_));
 sky130_fd_sc_hd__and2_2 _26861_ (.A(_16624_),
    .B(_16631_),
    .X(_16945_));
 sky130_fd_sc_hd__a21oi_2 _26862_ (.A1(_16622_),
    .A2(_16632_),
    .B1(_16945_),
    .Y(_16946_));
 sky130_fd_sc_hd__xor2_2 _26863_ (.A(_16944_),
    .B(_16946_),
    .X(_16948_));
 sky130_fd_sc_hd__xnor2_2 _26864_ (.A(_16930_),
    .B(_16948_),
    .Y(_16949_));
 sky130_fd_sc_hd__xor2_2 _26865_ (.A(_16906_),
    .B(_16949_),
    .X(_16950_));
 sky130_fd_sc_hd__xor2_2 _26866_ (.A(_16905_),
    .B(_16950_),
    .X(_16951_));
 sky130_fd_sc_hd__or2_2 _26867_ (.A(_16646_),
    .B(_16654_),
    .X(_16952_));
 sky130_fd_sc_hd__o21ai_2 _26868_ (.A1(_16652_),
    .A2(_16653_),
    .B1(_16952_),
    .Y(_16953_));
 sky130_fd_sc_hd__and2_2 _26869_ (.A(_16661_),
    .B(_16667_),
    .X(_16954_));
 sky130_fd_sc_hd__a21o_2 _26870_ (.A1(_16660_),
    .A2(_16668_),
    .B1(_16954_),
    .X(_16955_));
 sky130_fd_sc_hd__and4_2 _26871_ (.A(_13501_),
    .B(_13244_),
    .C(_14409_),
    .D(_14604_),
    .X(_16956_));
 sky130_fd_sc_hd__a22o_2 _26872_ (.A1(_14652_),
    .A2(_14410_),
    .B1(_14605_),
    .B2(_13501_),
    .X(_16957_));
 sky130_fd_sc_hd__and2b_2 _26873_ (.A_N(_16956_),
    .B(_16957_),
    .X(_16958_));
 sky130_fd_sc_hd__nor2_2 _26874_ (.A(_14343_),
    .B(_14948_),
    .Y(_16959_));
 sky130_fd_sc_hd__xnor2_2 _26875_ (.A(_16958_),
    .B(_16959_),
    .Y(_16960_));
 sky130_fd_sc_hd__nand2_2 _26876_ (.A(_13542_),
    .B(_13938_),
    .Y(_16961_));
 sky130_fd_sc_hd__xnor2_2 _26877_ (.A(_16647_),
    .B(_16961_),
    .Y(_16962_));
 sky130_fd_sc_hd__nand2_2 _26878_ (.A(_14648_),
    .B(_14391_),
    .Y(_16963_));
 sky130_fd_sc_hd__xnor2_2 _26879_ (.A(_16962_),
    .B(_16963_),
    .Y(_16964_));
 sky130_fd_sc_hd__o22a_2 _26880_ (.A1(_16275_),
    .A2(_16647_),
    .B1(_16648_),
    .B2(_16650_),
    .X(_16965_));
 sky130_fd_sc_hd__xnor2_2 _26881_ (.A(_16964_),
    .B(_16965_),
    .Y(_16966_));
 sky130_fd_sc_hd__xor2_2 _26882_ (.A(_16960_),
    .B(_16966_),
    .X(_16967_));
 sky130_fd_sc_hd__xnor2_2 _26883_ (.A(_16955_),
    .B(_16967_),
    .Y(_16969_));
 sky130_fd_sc_hd__xor2_2 _26884_ (.A(_16953_),
    .B(_16969_),
    .X(_16970_));
 sky130_fd_sc_hd__and2b_2 _26885_ (.A_N(_16665_),
    .B(_16666_),
    .X(_16971_));
 sky130_fd_sc_hd__a31o_2 _26886_ (.A1(_14637_),
    .A2(_16292_),
    .A3(_16663_),
    .B1(_16971_),
    .X(_16972_));
 sky130_fd_sc_hd__a21bo_2 _26887_ (.A1(_16670_),
    .A2(_16674_),
    .B1_N(_16672_),
    .X(_16973_));
 sky130_fd_sc_hd__nand2_2 _26888_ (.A(_12845_),
    .B(_14999_),
    .Y(_16974_));
 sky130_fd_sc_hd__and3_2 _26889_ (.A(_14634_),
    .B(_14994_),
    .C(_14996_),
    .X(_16975_));
 sky130_fd_sc_hd__xnor2_2 _26890_ (.A(_16974_),
    .B(_16975_),
    .Y(_16976_));
 sky130_fd_sc_hd__nor2_2 _26891_ (.A(_14641_),
    .B(_14988_),
    .Y(_16977_));
 sky130_fd_sc_hd__xnor2_2 _26892_ (.A(_16976_),
    .B(_16977_),
    .Y(_16978_));
 sky130_fd_sc_hd__xnor2_2 _26893_ (.A(_16973_),
    .B(_16978_),
    .Y(_16980_));
 sky130_fd_sc_hd__xnor2_2 _26894_ (.A(_16972_),
    .B(_16980_),
    .Y(_16981_));
 sky130_fd_sc_hd__and3_2 _26895_ (.A(_12242_),
    .B(_15900_),
    .C(_16671_),
    .X(_16982_));
 sky130_fd_sc_hd__nor2_2 _26896_ (.A(_13926_),
    .B(_16677_),
    .Y(_16983_));
 sky130_fd_sc_hd__a21o_2 _26897_ (.A1(_12242_),
    .A2(_15672_),
    .B1(_16983_),
    .X(_16984_));
 sky130_fd_sc_hd__and2b_2 _26898_ (.A_N(_16982_),
    .B(_16984_),
    .X(_16985_));
 sky130_fd_sc_hd__or3_2 _26899_ (.A(_14356_),
    .B(_15219_),
    .C(_15220_),
    .X(_16986_));
 sky130_fd_sc_hd__xnor2_2 _26900_ (.A(_16985_),
    .B(_16986_),
    .Y(_16987_));
 sky130_fd_sc_hd__buf_1 _26901_ (.A(_16689_),
    .X(_16988_));
 sky130_fd_sc_hd__and2_2 _26902_ (.A(iX[20]),
    .B(iX[52]),
    .X(_16989_));
 sky130_fd_sc_hd__nor2_2 _26903_ (.A(iX[20]),
    .B(iX[52]),
    .Y(_16991_));
 sky130_fd_sc_hd__or2_2 _26904_ (.A(_16989_),
    .B(_16991_),
    .X(_16992_));
 sky130_fd_sc_hd__buf_4 _26905_ (.A(_16992_),
    .X(_16993_));
 sky130_fd_sc_hd__nor4_2 _26906_ (.A(_15671_),
    .B(_15897_),
    .C(_16317_),
    .D(_16678_),
    .Y(_16994_));
 sky130_fd_sc_hd__and4bb_2 _26907_ (.A_N(_16317_),
    .B_N(_16678_),
    .C(_16315_),
    .D(_15894_),
    .X(_16995_));
 sky130_fd_sc_hd__o211a_2 _26908_ (.A1(iX[19]),
    .A2(iX[51]),
    .B1(iX[50]),
    .C1(iX[18]),
    .X(_16996_));
 sky130_fd_sc_hd__a211o_2 _26909_ (.A1(iX[19]),
    .A2(iX[51]),
    .B1(_16995_),
    .C1(_16996_),
    .X(_16997_));
 sky130_fd_sc_hd__a21oi_4 _26910_ (.A1(_15663_),
    .A2(_16994_),
    .B1(_16997_),
    .Y(_16998_));
 sky130_fd_sc_hd__xnor2_2 _26911_ (.A(_16993_),
    .B(_16998_),
    .Y(_16999_));
 sky130_fd_sc_hd__nor2_2 _26912_ (.A(_11575_),
    .B(_16999_),
    .Y(_17000_));
 sky130_fd_sc_hd__and3_2 _26913_ (.A(_11380_),
    .B(_16680_),
    .C(_17000_),
    .X(_17002_));
 sky130_fd_sc_hd__xor2_2 _26914_ (.A(_16993_),
    .B(_16998_),
    .X(_17003_));
 sky130_fd_sc_hd__a22o_2 _26915_ (.A1(_11583_),
    .A2(_16680_),
    .B1(_17003_),
    .B2(_11380_),
    .X(_17004_));
 sky130_fd_sc_hd__or4b_4 _26916_ (.A(_11793_),
    .B(_16988_),
    .C(_17002_),
    .D_N(_17004_),
    .X(_17005_));
 sky130_fd_sc_hd__buf_1 _26917_ (.A(_16682_),
    .X(_17006_));
 sky130_fd_sc_hd__buf_2 _26918_ (.A(_16686_),
    .X(_17007_));
 sky130_fd_sc_hd__or3b_2 _26919_ (.A(_11566_),
    .B(_17007_),
    .C_N(_17000_),
    .X(_17008_));
 sky130_fd_sc_hd__a22o_2 _26920_ (.A1(_15675_),
    .A2(_17006_),
    .B1(_17008_),
    .B2(_17004_),
    .X(_17009_));
 sky130_fd_sc_hd__a31o_2 _26921_ (.A1(_15675_),
    .A2(_15900_),
    .A3(_16683_),
    .B1(_16681_),
    .X(_17010_));
 sky130_fd_sc_hd__nand3_2 _26922_ (.A(_17005_),
    .B(_17009_),
    .C(_17010_),
    .Y(_17011_));
 sky130_fd_sc_hd__a21o_2 _26923_ (.A1(_17005_),
    .A2(_17009_),
    .B1(_17010_),
    .X(_17013_));
 sky130_fd_sc_hd__nand3_2 _26924_ (.A(_16987_),
    .B(_17011_),
    .C(_17013_),
    .Y(_17014_));
 sky130_fd_sc_hd__a21o_2 _26925_ (.A1(_17011_),
    .A2(_17013_),
    .B1(_16987_),
    .X(_17015_));
 sky130_fd_sc_hd__and3_2 _26926_ (.A(_16685_),
    .B(_16688_),
    .C(_16691_),
    .X(_17016_));
 sky130_fd_sc_hd__a31o_2 _26927_ (.A1(_16675_),
    .A2(_16676_),
    .A3(_16693_),
    .B1(_17016_),
    .X(_17017_));
 sky130_fd_sc_hd__and3_4 _26928_ (.A(_17014_),
    .B(_17015_),
    .C(_17017_),
    .X(_17018_));
 sky130_fd_sc_hd__a21oi_2 _26929_ (.A1(_17014_),
    .A2(_17015_),
    .B1(_17017_),
    .Y(_17019_));
 sky130_fd_sc_hd__or3_4 _26930_ (.A(_16981_),
    .B(_17018_),
    .C(_17019_),
    .X(_17020_));
 sky130_fd_sc_hd__o21ai_2 _26931_ (.A1(_17018_),
    .A2(_17019_),
    .B1(_16981_),
    .Y(_17021_));
 sky130_fd_sc_hd__o211a_2 _26932_ (.A1(_16698_),
    .A2(_16700_),
    .B1(_17020_),
    .C1(_17021_),
    .X(_17022_));
 sky130_fd_sc_hd__a211oi_2 _26933_ (.A1(_17020_),
    .A2(_17021_),
    .B1(_16698_),
    .C1(_16700_),
    .Y(_17024_));
 sky130_fd_sc_hd__or3_2 _26934_ (.A(_16970_),
    .B(_17022_),
    .C(_17024_),
    .X(_17025_));
 sky130_fd_sc_hd__o21ai_2 _26935_ (.A1(_17022_),
    .A2(_17024_),
    .B1(_16970_),
    .Y(_17026_));
 sky130_fd_sc_hd__nand2_2 _26936_ (.A(_17025_),
    .B(_17026_),
    .Y(_17027_));
 sky130_fd_sc_hd__nor2_2 _26937_ (.A(_16702_),
    .B(_16703_),
    .Y(_17028_));
 sky130_fd_sc_hd__a21oi_2 _26938_ (.A1(_16659_),
    .A2(_16704_),
    .B1(_17028_),
    .Y(_17029_));
 sky130_fd_sc_hd__xor2_2 _26939_ (.A(_17027_),
    .B(_17029_),
    .X(_17030_));
 sky130_fd_sc_hd__xnor2_2 _26940_ (.A(_16951_),
    .B(_17030_),
    .Y(_17031_));
 sky130_fd_sc_hd__nor2_2 _26941_ (.A(_16705_),
    .B(_16708_),
    .Y(_17032_));
 sky130_fd_sc_hd__nand2_2 _26942_ (.A(_16705_),
    .B(_16708_),
    .Y(_17033_));
 sky130_fd_sc_hd__o21a_2 _26943_ (.A1(_16638_),
    .A2(_17032_),
    .B1(_17033_),
    .X(_17035_));
 sky130_fd_sc_hd__nor2_2 _26944_ (.A(_17031_),
    .B(_17035_),
    .Y(_17036_));
 sky130_fd_sc_hd__nand2_2 _26945_ (.A(_17031_),
    .B(_17035_),
    .Y(_17037_));
 sky130_fd_sc_hd__and2b_2 _26946_ (.A_N(_17036_),
    .B(_17037_),
    .X(_17038_));
 sky130_fd_sc_hd__xnor2_2 _26947_ (.A(_16904_),
    .B(_17038_),
    .Y(_17039_));
 sky130_fd_sc_hd__or2b_2 _26948_ (.A(_16710_),
    .B_N(_16712_),
    .X(_17040_));
 sky130_fd_sc_hd__a21boi_2 _26949_ (.A1(_16601_),
    .A2(_16713_),
    .B1_N(_17040_),
    .Y(_17041_));
 sky130_fd_sc_hd__xor2_2 _26950_ (.A(_17039_),
    .B(_17041_),
    .X(_17042_));
 sky130_fd_sc_hd__xor2_2 _26951_ (.A(_16901_),
    .B(_17042_),
    .X(_17043_));
 sky130_fd_sc_hd__xnor2_2 _26952_ (.A(_16895_),
    .B(_17043_),
    .Y(_17044_));
 sky130_fd_sc_hd__xnor2_2 _26953_ (.A(_16900_),
    .B(_17044_),
    .Y(_17046_));
 sky130_fd_sc_hd__and2b_2 _26954_ (.A_N(_16582_),
    .B(_16583_),
    .X(_17047_));
 sky130_fd_sc_hd__and2_2 _26955_ (.A(_16584_),
    .B(_16586_),
    .X(_17048_));
 sky130_fd_sc_hd__nand3b_2 _26956_ (.A_N(_16581_),
    .B(_16551_),
    .C(_16550_),
    .Y(_17049_));
 sky130_fd_sc_hd__and3_2 _26957_ (.A(_16542_),
    .B(_16543_),
    .C(_16545_),
    .X(_17050_));
 sky130_fd_sc_hd__and2b_2 _26958_ (.A_N(_16503_),
    .B(_16502_),
    .X(_17051_));
 sky130_fd_sc_hd__or2b_2 _26959_ (.A(_16533_),
    .B_N(_16538_),
    .X(_17052_));
 sky130_fd_sc_hd__or2b_2 _26960_ (.A(_16532_),
    .B_N(_16539_),
    .X(_17053_));
 sky130_fd_sc_hd__and4_2 _26961_ (.A(iX[39]),
    .B(iX[40]),
    .C(iY[44]),
    .D(iY[45]),
    .X(_17054_));
 sky130_fd_sc_hd__a22oi_2 _26962_ (.A1(iX[40]),
    .A2(iY[44]),
    .B1(iY[45]),
    .B2(iX[39]),
    .Y(_17055_));
 sky130_fd_sc_hd__nor2_2 _26963_ (.A(_17054_),
    .B(_17055_),
    .Y(_17057_));
 sky130_fd_sc_hd__nand2_2 _26964_ (.A(iX[38]),
    .B(iY[46]),
    .Y(_17058_));
 sky130_fd_sc_hd__xnor2_2 _26965_ (.A(_17057_),
    .B(_17058_),
    .Y(_17059_));
 sky130_fd_sc_hd__and4_2 _26966_ (.A(iY[41]),
    .B(iX[42]),
    .C(iY[42]),
    .D(iX[43]),
    .X(_17060_));
 sky130_fd_sc_hd__a22oi_2 _26967_ (.A1(iX[42]),
    .A2(iY[42]),
    .B1(iX[43]),
    .B2(iY[41]),
    .Y(_17061_));
 sky130_fd_sc_hd__nor2_2 _26968_ (.A(_17060_),
    .B(_17061_),
    .Y(_17062_));
 sky130_fd_sc_hd__nand2_2 _26969_ (.A(iX[41]),
    .B(iY[43]),
    .Y(_17063_));
 sky130_fd_sc_hd__xnor2_2 _26970_ (.A(_17062_),
    .B(_17063_),
    .Y(_17064_));
 sky130_fd_sc_hd__o21ba_2 _26971_ (.A1(_16499_),
    .A2(_16501_),
    .B1_N(_16498_),
    .X(_17065_));
 sky130_fd_sc_hd__xnor2_2 _26972_ (.A(_17064_),
    .B(_17065_),
    .Y(_17066_));
 sky130_fd_sc_hd__and2_2 _26973_ (.A(_17059_),
    .B(_17066_),
    .X(_17068_));
 sky130_fd_sc_hd__nor2_2 _26974_ (.A(_17059_),
    .B(_17066_),
    .Y(_17069_));
 sky130_fd_sc_hd__or2_2 _26975_ (.A(_17068_),
    .B(_17069_),
    .X(_17070_));
 sky130_fd_sc_hd__a21o_2 _26976_ (.A1(_17052_),
    .A2(_17053_),
    .B1(_17070_),
    .X(_17071_));
 sky130_fd_sc_hd__nand3_2 _26977_ (.A(_17052_),
    .B(_17053_),
    .C(_17070_),
    .Y(_17072_));
 sky130_fd_sc_hd__o211ai_2 _26978_ (.A1(_17051_),
    .A2(_16505_),
    .B1(_17071_),
    .C1(_17072_),
    .Y(_17073_));
 sky130_fd_sc_hd__a211o_2 _26979_ (.A1(_17071_),
    .A2(_17072_),
    .B1(_17051_),
    .C1(_16505_),
    .X(_17074_));
 sky130_fd_sc_hd__or2b_2 _26980_ (.A(_16521_),
    .B_N(_16520_),
    .X(_17075_));
 sky130_fd_sc_hd__nand2_2 _26981_ (.A(_16522_),
    .B(_16527_),
    .Y(_17076_));
 sky130_fd_sc_hd__and4_2 _26982_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[49]),
    .D(iX[50]),
    .X(_17077_));
 sky130_fd_sc_hd__a22oi_2 _26983_ (.A1(iY[35]),
    .A2(iX[49]),
    .B1(iX[50]),
    .B2(iY[34]),
    .Y(_17079_));
 sky130_fd_sc_hd__nor2_2 _26984_ (.A(_17077_),
    .B(_17079_),
    .Y(_17080_));
 sky130_fd_sc_hd__nand2_2 _26985_ (.A(iY[33]),
    .B(iX[51]),
    .Y(_17081_));
 sky130_fd_sc_hd__xnor2_2 _26986_ (.A(_17080_),
    .B(_17081_),
    .Y(_17082_));
 sky130_fd_sc_hd__o21ba_2 _26987_ (.A1(_16516_),
    .A2(_16518_),
    .B1_N(_16515_),
    .X(_17083_));
 sky130_fd_sc_hd__xnor2_2 _26988_ (.A(_17082_),
    .B(_17083_),
    .Y(_17084_));
 sky130_fd_sc_hd__and4_2 _26989_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[48]),
    .D(iX[52]),
    .X(_17085_));
 sky130_fd_sc_hd__a22oi_2 _26990_ (.A1(iY[36]),
    .A2(iX[48]),
    .B1(iX[52]),
    .B2(iY[32]),
    .Y(_17086_));
 sky130_fd_sc_hd__nor2_2 _26991_ (.A(_17085_),
    .B(_17086_),
    .Y(_17087_));
 sky130_fd_sc_hd__nand2_2 _26992_ (.A(iY[37]),
    .B(iX[47]),
    .Y(_17088_));
 sky130_fd_sc_hd__xnor2_2 _26993_ (.A(_17087_),
    .B(_17088_),
    .Y(_17090_));
 sky130_fd_sc_hd__xnor2_2 _26994_ (.A(_17084_),
    .B(_17090_),
    .Y(_17091_));
 sky130_fd_sc_hd__a21o_2 _26995_ (.A1(_17075_),
    .A2(_17076_),
    .B1(_17091_),
    .X(_17092_));
 sky130_fd_sc_hd__nand3_2 _26996_ (.A(_17075_),
    .B(_17076_),
    .C(_17091_),
    .Y(_17093_));
 sky130_fd_sc_hd__o21ba_2 _26997_ (.A1(_16535_),
    .A2(_16537_),
    .B1_N(_16534_),
    .X(_17094_));
 sky130_fd_sc_hd__o21ba_2 _26998_ (.A1(_16524_),
    .A2(_16526_),
    .B1_N(_16523_),
    .X(_17095_));
 sky130_fd_sc_hd__and4_2 _26999_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[45]),
    .D(iX[46]),
    .X(_17096_));
 sky130_fd_sc_hd__a22oi_2 _27000_ (.A1(iY[39]),
    .A2(iX[45]),
    .B1(iX[46]),
    .B2(iY[38]),
    .Y(_17097_));
 sky130_fd_sc_hd__nor2_2 _27001_ (.A(_17096_),
    .B(_17097_),
    .Y(_17098_));
 sky130_fd_sc_hd__nand2_2 _27002_ (.A(iY[40]),
    .B(iX[44]),
    .Y(_17099_));
 sky130_fd_sc_hd__xnor2_2 _27003_ (.A(_17098_),
    .B(_17099_),
    .Y(_17101_));
 sky130_fd_sc_hd__xnor2_2 _27004_ (.A(_17095_),
    .B(_17101_),
    .Y(_17102_));
 sky130_fd_sc_hd__xnor2_2 _27005_ (.A(_17094_),
    .B(_17102_),
    .Y(_17103_));
 sky130_fd_sc_hd__nand3_2 _27006_ (.A(_17092_),
    .B(_17093_),
    .C(_17103_),
    .Y(_17104_));
 sky130_fd_sc_hd__a21o_2 _27007_ (.A1(_17092_),
    .A2(_17093_),
    .B1(_17103_),
    .X(_17105_));
 sky130_fd_sc_hd__nand2_2 _27008_ (.A(_17104_),
    .B(_17105_),
    .Y(_17106_));
 sky130_fd_sc_hd__nand2_2 _27009_ (.A(_16529_),
    .B(_16542_),
    .Y(_17107_));
 sky130_fd_sc_hd__xnor2_2 _27010_ (.A(_17106_),
    .B(_17107_),
    .Y(_17108_));
 sky130_fd_sc_hd__a21o_2 _27011_ (.A1(_17073_),
    .A2(_17074_),
    .B1(_17108_),
    .X(_17109_));
 sky130_fd_sc_hd__and3_2 _27012_ (.A(_17108_),
    .B(_17073_),
    .C(_17074_),
    .X(_17110_));
 sky130_fd_sc_hd__inv_2 _27013_ (.A(_17110_),
    .Y(_17112_));
 sky130_fd_sc_hd__o211a_2 _27014_ (.A1(_17050_),
    .A2(_16548_),
    .B1(_17109_),
    .C1(_17112_),
    .X(_17113_));
 sky130_fd_sc_hd__a211oi_2 _27015_ (.A1(_17109_),
    .A2(_17112_),
    .B1(_17050_),
    .C1(_16548_),
    .Y(_17114_));
 sky130_fd_sc_hd__and4_2 _27016_ (.A(iX[33]),
    .B(iX[34]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_17115_));
 sky130_fd_sc_hd__a22oi_2 _27017_ (.A1(iX[34]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[33]),
    .Y(_17116_));
 sky130_fd_sc_hd__nor2_2 _27018_ (.A(_17115_),
    .B(_17116_),
    .Y(_17117_));
 sky130_fd_sc_hd__nand2_2 _27019_ (.A(iX[32]),
    .B(iY[52]),
    .Y(_17118_));
 sky130_fd_sc_hd__xnor2_2 _27020_ (.A(_17117_),
    .B(_17118_),
    .Y(_17119_));
 sky130_fd_sc_hd__and2_2 _27021_ (.A(_16557_),
    .B(_17119_),
    .X(_17120_));
 sky130_fd_sc_hd__nor2_2 _27022_ (.A(_16557_),
    .B(_17119_),
    .Y(_17121_));
 sky130_fd_sc_hd__or2_2 _27023_ (.A(_17120_),
    .B(_17121_),
    .X(_17123_));
 sky130_fd_sc_hd__or3_2 _27024_ (.A(_16560_),
    .B(_16565_),
    .C(_16566_),
    .X(_17124_));
 sky130_fd_sc_hd__nand2_2 _27025_ (.A(_16559_),
    .B(_16568_),
    .Y(_17125_));
 sky130_fd_sc_hd__o21ba_2 _27026_ (.A1(_16493_),
    .A2(_16495_),
    .B1_N(_16492_),
    .X(_17126_));
 sky130_fd_sc_hd__and4_2 _27027_ (.A(iX[36]),
    .B(iX[37]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_17127_));
 sky130_fd_sc_hd__a22oi_2 _27028_ (.A1(iX[37]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[36]),
    .Y(_17128_));
 sky130_fd_sc_hd__nand2_2 _27029_ (.A(iX[35]),
    .B(iY[49]),
    .Y(_17129_));
 sky130_fd_sc_hd__o21a_2 _27030_ (.A1(_17127_),
    .A2(_17128_),
    .B1(_17129_),
    .X(_17130_));
 sky130_fd_sc_hd__nor3_2 _27031_ (.A(_17127_),
    .B(_17128_),
    .C(_17129_),
    .Y(_17131_));
 sky130_fd_sc_hd__nor2_2 _27032_ (.A(_17130_),
    .B(_17131_),
    .Y(_17132_));
 sky130_fd_sc_hd__xnor2_2 _27033_ (.A(_17126_),
    .B(_17132_),
    .Y(_17134_));
 sky130_fd_sc_hd__o21ai_2 _27034_ (.A1(_16561_),
    .A2(_16566_),
    .B1(_17134_),
    .Y(_17135_));
 sky130_fd_sc_hd__or3_2 _27035_ (.A(_16561_),
    .B(_16566_),
    .C(_17134_),
    .X(_17136_));
 sky130_fd_sc_hd__nand2_2 _27036_ (.A(_17135_),
    .B(_17136_),
    .Y(_17137_));
 sky130_fd_sc_hd__a21oi_2 _27037_ (.A1(_17124_),
    .A2(_17125_),
    .B1(_17137_),
    .Y(_17138_));
 sky130_fd_sc_hd__and3_2 _27038_ (.A(_17124_),
    .B(_17125_),
    .C(_17137_),
    .X(_17139_));
 sky130_fd_sc_hd__or3_2 _27039_ (.A(_17123_),
    .B(_17138_),
    .C(_17139_),
    .X(_17140_));
 sky130_fd_sc_hd__o21ai_2 _27040_ (.A1(_17138_),
    .A2(_17139_),
    .B1(_17123_),
    .Y(_17141_));
 sky130_fd_sc_hd__nand2_2 _27041_ (.A(_17140_),
    .B(_17141_),
    .Y(_17142_));
 sky130_fd_sc_hd__a21oi_2 _27042_ (.A1(_16509_),
    .A2(_16511_),
    .B1(_17142_),
    .Y(_17143_));
 sky130_fd_sc_hd__and3_2 _27043_ (.A(_16509_),
    .B(_16511_),
    .C(_17142_),
    .X(_17145_));
 sky130_fd_sc_hd__a211oi_2 _27044_ (.A1(_16570_),
    .A2(_16573_),
    .B1(_17143_),
    .C1(_17145_),
    .Y(_17146_));
 sky130_fd_sc_hd__o211a_2 _27045_ (.A1(_17143_),
    .A2(_17145_),
    .B1(_16570_),
    .C1(_16573_),
    .X(_17147_));
 sky130_fd_sc_hd__nor4_2 _27046_ (.A(_17113_),
    .B(_17114_),
    .C(_17146_),
    .D(_17147_),
    .Y(_17148_));
 sky130_fd_sc_hd__o22a_2 _27047_ (.A1(_17113_),
    .A2(_17114_),
    .B1(_17146_),
    .B2(_17147_),
    .X(_17149_));
 sky130_fd_sc_hd__a211oi_2 _27048_ (.A1(_16550_),
    .A2(_17049_),
    .B1(_17148_),
    .C1(_17149_),
    .Y(_17150_));
 sky130_fd_sc_hd__o211a_2 _27049_ (.A1(_17148_),
    .A2(_17149_),
    .B1(_16550_),
    .C1(_17049_),
    .X(_17151_));
 sky130_fd_sc_hd__nor2_2 _27050_ (.A(_16576_),
    .B(_16579_),
    .Y(_17152_));
 sky130_fd_sc_hd__or3_2 _27051_ (.A(_17150_),
    .B(_17151_),
    .C(_17152_),
    .X(_17153_));
 sky130_fd_sc_hd__o21ai_2 _27052_ (.A1(_17150_),
    .A2(_17151_),
    .B1(_17152_),
    .Y(_17154_));
 sky130_fd_sc_hd__nand2_2 _27053_ (.A(_17153_),
    .B(_17154_),
    .Y(_17156_));
 sky130_fd_sc_hd__o21ba_2 _27054_ (.A1(_17047_),
    .A2(_17048_),
    .B1_N(_17156_),
    .X(_17157_));
 sky130_fd_sc_hd__nor3b_2 _27055_ (.A(_17047_),
    .B(_17048_),
    .C_N(_17156_),
    .Y(_17158_));
 sky130_fd_sc_hd__or3_2 _27056_ (.A(_16588_),
    .B(_17157_),
    .C(_17158_),
    .X(_17159_));
 sky130_fd_sc_hd__o21ai_2 _27057_ (.A1(_17157_),
    .A2(_17158_),
    .B1(_16588_),
    .Y(_17160_));
 sky130_fd_sc_hd__and2_2 _27058_ (.A(_17159_),
    .B(_17160_),
    .X(_17161_));
 sky130_fd_sc_hd__xor2_2 _27059_ (.A(_16590_),
    .B(_17161_),
    .X(_17162_));
 sky130_fd_sc_hd__a21oi_2 _27060_ (.A1(_16028_),
    .A2(_16032_),
    .B1(_16029_),
    .Y(_17163_));
 sky130_fd_sc_hd__and2b_2 _27061_ (.A_N(_16593_),
    .B(_16458_),
    .X(_17164_));
 sky130_fd_sc_hd__a311oi_2 _27062_ (.A1(_15713_),
    .A2(_15806_),
    .A3(_16026_),
    .B1(_16592_),
    .C1(_17164_),
    .Y(_17165_));
 sky130_fd_sc_hd__o21ba_2 _27063_ (.A1(_16457_),
    .A2(_16593_),
    .B1_N(_16592_),
    .X(_17167_));
 sky130_fd_sc_hd__a21o_2 _27064_ (.A1(_17163_),
    .A2(_17165_),
    .B1(_17167_),
    .X(_17168_));
 sky130_fd_sc_hd__nor2_2 _27065_ (.A(_17162_),
    .B(_17168_),
    .Y(_17169_));
 sky130_fd_sc_hd__and2_2 _27066_ (.A(_17162_),
    .B(_17168_),
    .X(_17170_));
 sky130_fd_sc_hd__nor2_2 _27067_ (.A(_17169_),
    .B(_17170_),
    .Y(_17171_));
 sky130_fd_sc_hd__nand2_2 _27068_ (.A(_17046_),
    .B(_17171_),
    .Y(_17172_));
 sky130_fd_sc_hd__or2_2 _27069_ (.A(_17046_),
    .B(_17171_),
    .X(_17173_));
 sky130_fd_sc_hd__nand2_2 _27070_ (.A(_17172_),
    .B(_17173_),
    .Y(_17174_));
 sky130_fd_sc_hd__xnor2_2 _27071_ (.A(oO[20]),
    .B(_17174_),
    .Y(_17175_));
 sky130_fd_sc_hd__inv_2 _27072_ (.A(_16597_),
    .Y(_17176_));
 sky130_fd_sc_hd__nor2_2 _27073_ (.A(_17176_),
    .B(_16722_),
    .Y(_17178_));
 sky130_fd_sc_hd__a21oi_2 _27074_ (.A1(_03114_),
    .A2(_16723_),
    .B1(_17178_),
    .Y(_17179_));
 sky130_fd_sc_hd__xnor2_2 _27075_ (.A(_17175_),
    .B(_17179_),
    .Y(_17180_));
 sky130_fd_sc_hd__a21oi_2 _27076_ (.A1(_16891_),
    .A2(_16732_),
    .B1(_17180_),
    .Y(_17181_));
 sky130_fd_sc_hd__and3_2 _27077_ (.A(_16891_),
    .B(_16732_),
    .C(_17180_),
    .X(_17182_));
 sky130_fd_sc_hd__nor2_2 _27078_ (.A(_17181_),
    .B(_17182_),
    .Y(_17183_));
 sky130_fd_sc_hd__xor2_2 _27079_ (.A(_16890_),
    .B(_17183_),
    .X(_17184_));
 sky130_fd_sc_hd__and2b_2 _27080_ (.A_N(_16810_),
    .B(_16478_),
    .X(_17185_));
 sky130_fd_sc_hd__nor2_2 _27081_ (.A(_16811_),
    .B(_17185_),
    .Y(_17186_));
 sky130_fd_sc_hd__and2_2 _27082_ (.A(_16482_),
    .B(_17186_),
    .X(_17187_));
 sky130_fd_sc_hd__nand2_2 _27083_ (.A(_16480_),
    .B(_16812_),
    .Y(_17189_));
 sky130_fd_sc_hd__a22oi_2 _27084_ (.A1(_16481_),
    .A2(_17187_),
    .B1(_17189_),
    .B2(_17186_),
    .Y(_17190_));
 sky130_fd_sc_hd__xnor2_2 _27085_ (.A(_17184_),
    .B(_17190_),
    .Y(oO[52]));
 sky130_fd_sc_hd__and2b_2 _27086_ (.A_N(_16886_),
    .B(_16885_),
    .X(_17191_));
 sky130_fd_sc_hd__or2_2 _27087_ (.A(_17191_),
    .B(_16888_),
    .X(_17192_));
 sky130_fd_sc_hd__or2b_2 _27088_ (.A(_16883_),
    .B_N(_16884_),
    .X(_17193_));
 sky130_fd_sc_hd__a22o_2 _27089_ (.A1(iY[23]),
    .A2(iX[30]),
    .B1(iX[31]),
    .B2(iY[22]),
    .X(_17194_));
 sky130_fd_sc_hd__and3_2 _27090_ (.A(iY[23]),
    .B(iX[31]),
    .C(_16736_),
    .X(_17195_));
 sky130_fd_sc_hd__inv_2 _27091_ (.A(_17195_),
    .Y(_17196_));
 sky130_fd_sc_hd__o21ba_2 _27092_ (.A1(_16832_),
    .A2(_16834_),
    .B1_N(_16831_),
    .X(_17197_));
 sky130_fd_sc_hd__a31o_2 _27093_ (.A1(iY[23]),
    .A2(iX[29]),
    .A3(_16820_),
    .B1(_16819_),
    .X(_17199_));
 sky130_fd_sc_hd__and4_2 _27094_ (.A(iY[24]),
    .B(iY[25]),
    .C(iX[28]),
    .D(iX[29]),
    .X(_17200_));
 sky130_fd_sc_hd__a22oi_2 _27095_ (.A1(iY[25]),
    .A2(iX[28]),
    .B1(iX[29]),
    .B2(iY[24]),
    .Y(_17201_));
 sky130_fd_sc_hd__nor2_2 _27096_ (.A(_17200_),
    .B(_17201_),
    .Y(_17202_));
 sky130_fd_sc_hd__nand2_2 _27097_ (.A(iY[26]),
    .B(iX[27]),
    .Y(_17203_));
 sky130_fd_sc_hd__xnor2_2 _27098_ (.A(_17202_),
    .B(_17203_),
    .Y(_17204_));
 sky130_fd_sc_hd__nand2_2 _27099_ (.A(_17199_),
    .B(_17204_),
    .Y(_17205_));
 sky130_fd_sc_hd__or2_2 _27100_ (.A(_17199_),
    .B(_17204_),
    .X(_17206_));
 sky130_fd_sc_hd__and2_2 _27101_ (.A(_17205_),
    .B(_17206_),
    .X(_17207_));
 sky130_fd_sc_hd__or2b_2 _27102_ (.A(_17197_),
    .B_N(_17207_),
    .X(_17208_));
 sky130_fd_sc_hd__or2b_2 _27103_ (.A(_17207_),
    .B_N(_17197_),
    .X(_17210_));
 sky130_fd_sc_hd__nand2_2 _27104_ (.A(_17208_),
    .B(_17210_),
    .Y(_17211_));
 sky130_fd_sc_hd__o21ba_2 _27105_ (.A1(_16830_),
    .A2(_16838_),
    .B1_N(_16836_),
    .X(_17212_));
 sky130_fd_sc_hd__or2_2 _27106_ (.A(_17211_),
    .B(_17212_),
    .X(_17213_));
 sky130_fd_sc_hd__nand2_2 _27107_ (.A(_17211_),
    .B(_17212_),
    .Y(_17214_));
 sky130_fd_sc_hd__nand2_2 _27108_ (.A(_17213_),
    .B(_17214_),
    .Y(_17215_));
 sky130_fd_sc_hd__inv_2 _27109_ (.A(_16829_),
    .Y(_17216_));
 sky130_fd_sc_hd__a21oi_2 _27110_ (.A1(_17216_),
    .A2(_16840_),
    .B1(_16842_),
    .Y(_17217_));
 sky130_fd_sc_hd__or2_2 _27111_ (.A(_17215_),
    .B(_17217_),
    .X(_17218_));
 sky130_fd_sc_hd__nand2_2 _27112_ (.A(_17215_),
    .B(_17217_),
    .Y(_17219_));
 sky130_fd_sc_hd__and2_2 _27113_ (.A(_17218_),
    .B(_17219_),
    .X(_17221_));
 sky130_fd_sc_hd__or2b_2 _27114_ (.A(_16854_),
    .B_N(_16853_),
    .X(_17222_));
 sky130_fd_sc_hd__and4_2 _27115_ (.A(iX[25]),
    .B(iX[26]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_17223_));
 sky130_fd_sc_hd__a22oi_2 _27116_ (.A1(iX[26]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[25]),
    .Y(_17224_));
 sky130_fd_sc_hd__nor2_2 _27117_ (.A(_17223_),
    .B(_17224_),
    .Y(_17225_));
 sky130_fd_sc_hd__nand2_2 _27118_ (.A(iX[24]),
    .B(iY[29]),
    .Y(_17226_));
 sky130_fd_sc_hd__xnor2_2 _27119_ (.A(_17225_),
    .B(_17226_),
    .Y(_17227_));
 sky130_fd_sc_hd__o21ba_2 _27120_ (.A1(_16850_),
    .A2(_16852_),
    .B1_N(_16849_),
    .X(_17228_));
 sky130_fd_sc_hd__xnor2_2 _27121_ (.A(_17227_),
    .B(_17228_),
    .Y(_17229_));
 sky130_fd_sc_hd__nand3_2 _27122_ (.A(iX[23]),
    .B(iY[30]),
    .C(_17229_),
    .Y(_17230_));
 sky130_fd_sc_hd__a21o_2 _27123_ (.A1(iX[23]),
    .A2(iY[30]),
    .B1(_17229_),
    .X(_17232_));
 sky130_fd_sc_hd__nand2_2 _27124_ (.A(_17230_),
    .B(_17232_),
    .Y(_17233_));
 sky130_fd_sc_hd__a21oi_2 _27125_ (.A1(_17222_),
    .A2(_16856_),
    .B1(_17233_),
    .Y(_17234_));
 sky130_fd_sc_hd__and3_2 _27126_ (.A(_17222_),
    .B(_16856_),
    .C(_17233_),
    .X(_17235_));
 sky130_fd_sc_hd__nor2_2 _27127_ (.A(_17234_),
    .B(_17235_),
    .Y(_17236_));
 sky130_fd_sc_hd__nand2_2 _27128_ (.A(iX[22]),
    .B(iY[31]),
    .Y(_17237_));
 sky130_fd_sc_hd__xnor2_2 _27129_ (.A(_17236_),
    .B(_17237_),
    .Y(_17238_));
 sky130_fd_sc_hd__nand2_2 _27130_ (.A(_17221_),
    .B(_17238_),
    .Y(_17239_));
 sky130_fd_sc_hd__or2_2 _27131_ (.A(_17221_),
    .B(_17238_),
    .X(_17240_));
 sky130_fd_sc_hd__and2_2 _27132_ (.A(_17239_),
    .B(_17240_),
    .X(_17241_));
 sky130_fd_sc_hd__nor2_2 _27133_ (.A(_16844_),
    .B(_16865_),
    .Y(_17243_));
 sky130_fd_sc_hd__xnor2_2 _27134_ (.A(_17241_),
    .B(_17243_),
    .Y(_17244_));
 sky130_fd_sc_hd__and3_2 _27135_ (.A(_17194_),
    .B(_17196_),
    .C(_17244_),
    .X(_17245_));
 sky130_fd_sc_hd__a21oi_2 _27136_ (.A1(_17194_),
    .A2(_17196_),
    .B1(_17244_),
    .Y(_17246_));
 sky130_fd_sc_hd__nor2_2 _27137_ (.A(_17245_),
    .B(_17246_),
    .Y(_17247_));
 sky130_fd_sc_hd__xnor2_2 _27138_ (.A(_16871_),
    .B(_17247_),
    .Y(_17248_));
 sky130_fd_sc_hd__xnor2_2 _27139_ (.A(_16867_),
    .B(_17248_),
    .Y(_17249_));
 sky130_fd_sc_hd__a21oi_2 _27140_ (.A1(_16874_),
    .A2(_16877_),
    .B1(_17249_),
    .Y(_17250_));
 sky130_fd_sc_hd__nand3_2 _27141_ (.A(_16874_),
    .B(_16877_),
    .C(_17249_),
    .Y(_17251_));
 sky130_fd_sc_hd__and2b_2 _27142_ (.A_N(_17250_),
    .B(_17251_),
    .X(_17252_));
 sky130_fd_sc_hd__a31o_2 _27143_ (.A1(iX[21]),
    .A2(iY[31]),
    .A3(_16862_),
    .B1(_16860_),
    .X(_17254_));
 sky130_fd_sc_hd__xnor2_2 _27144_ (.A(_17252_),
    .B(_17254_),
    .Y(_17255_));
 sky130_fd_sc_hd__a21oi_2 _27145_ (.A1(_16880_),
    .A2(_17193_),
    .B1(_17255_),
    .Y(_17256_));
 sky130_fd_sc_hd__and3_2 _27146_ (.A(_16880_),
    .B(_17193_),
    .C(_17255_),
    .X(_17257_));
 sky130_fd_sc_hd__nor2_2 _27147_ (.A(_17256_),
    .B(_17257_),
    .Y(_17258_));
 sky130_fd_sc_hd__xnor2_2 _27148_ (.A(_17192_),
    .B(_17258_),
    .Y(_17259_));
 sky130_fd_sc_hd__and2b_2 _27149_ (.A_N(_16590_),
    .B(_17161_),
    .X(_17260_));
 sky130_fd_sc_hd__and3_2 _27150_ (.A(_17104_),
    .B(_17105_),
    .C(_17107_),
    .X(_17261_));
 sky130_fd_sc_hd__and2b_2 _27151_ (.A_N(_17065_),
    .B(_17064_),
    .X(_17262_));
 sky130_fd_sc_hd__or2b_2 _27152_ (.A(_17095_),
    .B_N(_17101_),
    .X(_17263_));
 sky130_fd_sc_hd__or2b_2 _27153_ (.A(_17094_),
    .B_N(_17102_),
    .X(_17265_));
 sky130_fd_sc_hd__and4_2 _27154_ (.A(iX[40]),
    .B(iX[41]),
    .C(iY[44]),
    .D(iY[45]),
    .X(_17266_));
 sky130_fd_sc_hd__a22oi_2 _27155_ (.A1(iX[41]),
    .A2(iY[44]),
    .B1(iY[45]),
    .B2(iX[40]),
    .Y(_17267_));
 sky130_fd_sc_hd__nor2_2 _27156_ (.A(_17266_),
    .B(_17267_),
    .Y(_17268_));
 sky130_fd_sc_hd__nand2_2 _27157_ (.A(iX[39]),
    .B(iY[46]),
    .Y(_17269_));
 sky130_fd_sc_hd__xnor2_2 _27158_ (.A(_17268_),
    .B(_17269_),
    .Y(_17270_));
 sky130_fd_sc_hd__and4_2 _27159_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[43]),
    .D(iX[44]),
    .X(_17271_));
 sky130_fd_sc_hd__a22oi_2 _27160_ (.A1(iY[42]),
    .A2(iX[43]),
    .B1(iX[44]),
    .B2(iY[41]),
    .Y(_17272_));
 sky130_fd_sc_hd__nor2_2 _27161_ (.A(_17271_),
    .B(_17272_),
    .Y(_17273_));
 sky130_fd_sc_hd__nand2_2 _27162_ (.A(iX[42]),
    .B(iY[43]),
    .Y(_17274_));
 sky130_fd_sc_hd__xnor2_2 _27163_ (.A(_17273_),
    .B(_17274_),
    .Y(_17276_));
 sky130_fd_sc_hd__o21ba_2 _27164_ (.A1(_17061_),
    .A2(_17063_),
    .B1_N(_17060_),
    .X(_17277_));
 sky130_fd_sc_hd__xnor2_2 _27165_ (.A(_17276_),
    .B(_17277_),
    .Y(_17278_));
 sky130_fd_sc_hd__xnor2_2 _27166_ (.A(_17270_),
    .B(_17278_),
    .Y(_17279_));
 sky130_fd_sc_hd__a21o_2 _27167_ (.A1(_17263_),
    .A2(_17265_),
    .B1(_17279_),
    .X(_17280_));
 sky130_fd_sc_hd__nand3_2 _27168_ (.A(_17263_),
    .B(_17265_),
    .C(_17279_),
    .Y(_17281_));
 sky130_fd_sc_hd__o211ai_2 _27169_ (.A1(_17262_),
    .A2(_17068_),
    .B1(_17280_),
    .C1(_17281_),
    .Y(_17282_));
 sky130_fd_sc_hd__a211o_2 _27170_ (.A1(_17280_),
    .A2(_17281_),
    .B1(_17262_),
    .C1(_17068_),
    .X(_17283_));
 sky130_fd_sc_hd__or2b_2 _27171_ (.A(_17083_),
    .B_N(_17082_),
    .X(_17284_));
 sky130_fd_sc_hd__nand2_2 _27172_ (.A(_17084_),
    .B(_17090_),
    .Y(_17285_));
 sky130_fd_sc_hd__and4_2 _27173_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[50]),
    .D(iX[51]),
    .X(_17287_));
 sky130_fd_sc_hd__a22oi_2 _27174_ (.A1(iY[35]),
    .A2(iX[50]),
    .B1(iX[51]),
    .B2(iY[34]),
    .Y(_17288_));
 sky130_fd_sc_hd__nor2_2 _27175_ (.A(_17287_),
    .B(_17288_),
    .Y(_17289_));
 sky130_fd_sc_hd__nand2_2 _27176_ (.A(iY[33]),
    .B(iX[52]),
    .Y(_17290_));
 sky130_fd_sc_hd__xnor2_2 _27177_ (.A(_17289_),
    .B(_17290_),
    .Y(_17291_));
 sky130_fd_sc_hd__o21ba_2 _27178_ (.A1(_17079_),
    .A2(_17081_),
    .B1_N(_17077_),
    .X(_17292_));
 sky130_fd_sc_hd__xnor2_2 _27179_ (.A(_17291_),
    .B(_17292_),
    .Y(_17293_));
 sky130_fd_sc_hd__and4_2 _27180_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[49]),
    .D(iX[53]),
    .X(_17294_));
 sky130_fd_sc_hd__a22oi_2 _27181_ (.A1(iY[36]),
    .A2(iX[49]),
    .B1(iX[53]),
    .B2(iY[32]),
    .Y(_17295_));
 sky130_fd_sc_hd__nor2_2 _27182_ (.A(_17294_),
    .B(_17295_),
    .Y(_17296_));
 sky130_fd_sc_hd__nand2_2 _27183_ (.A(iY[37]),
    .B(iX[48]),
    .Y(_17298_));
 sky130_fd_sc_hd__xnor2_2 _27184_ (.A(_17296_),
    .B(_17298_),
    .Y(_17299_));
 sky130_fd_sc_hd__xnor2_2 _27185_ (.A(_17293_),
    .B(_17299_),
    .Y(_17300_));
 sky130_fd_sc_hd__a21o_2 _27186_ (.A1(_17284_),
    .A2(_17285_),
    .B1(_17300_),
    .X(_17301_));
 sky130_fd_sc_hd__nand3_2 _27187_ (.A(_17284_),
    .B(_17285_),
    .C(_17300_),
    .Y(_17302_));
 sky130_fd_sc_hd__o21ba_2 _27188_ (.A1(_17097_),
    .A2(_17099_),
    .B1_N(_17096_),
    .X(_17303_));
 sky130_fd_sc_hd__o21ba_2 _27189_ (.A1(_17086_),
    .A2(_17088_),
    .B1_N(_17085_),
    .X(_17304_));
 sky130_fd_sc_hd__and4_2 _27190_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[46]),
    .D(iX[47]),
    .X(_17305_));
 sky130_fd_sc_hd__a22oi_2 _27191_ (.A1(iY[39]),
    .A2(iX[46]),
    .B1(iX[47]),
    .B2(iY[38]),
    .Y(_17306_));
 sky130_fd_sc_hd__nor2_2 _27192_ (.A(_17305_),
    .B(_17306_),
    .Y(_17307_));
 sky130_fd_sc_hd__nand2_2 _27193_ (.A(iY[40]),
    .B(iX[45]),
    .Y(_17309_));
 sky130_fd_sc_hd__xnor2_2 _27194_ (.A(_17307_),
    .B(_17309_),
    .Y(_17310_));
 sky130_fd_sc_hd__xnor2_2 _27195_ (.A(_17304_),
    .B(_17310_),
    .Y(_17311_));
 sky130_fd_sc_hd__xnor2_2 _27196_ (.A(_17303_),
    .B(_17311_),
    .Y(_17312_));
 sky130_fd_sc_hd__nand3_2 _27197_ (.A(_17301_),
    .B(_17302_),
    .C(_17312_),
    .Y(_17313_));
 sky130_fd_sc_hd__a21o_2 _27198_ (.A1(_17301_),
    .A2(_17302_),
    .B1(_17312_),
    .X(_17314_));
 sky130_fd_sc_hd__nand2_2 _27199_ (.A(_17313_),
    .B(_17314_),
    .Y(_17315_));
 sky130_fd_sc_hd__nand2_2 _27200_ (.A(_17092_),
    .B(_17104_),
    .Y(_17316_));
 sky130_fd_sc_hd__xnor2_2 _27201_ (.A(_17315_),
    .B(_17316_),
    .Y(_17317_));
 sky130_fd_sc_hd__a21o_2 _27202_ (.A1(_17282_),
    .A2(_17283_),
    .B1(_17317_),
    .X(_17318_));
 sky130_fd_sc_hd__and3_2 _27203_ (.A(_17317_),
    .B(_17282_),
    .C(_17283_),
    .X(_17320_));
 sky130_fd_sc_hd__inv_2 _27204_ (.A(_17320_),
    .Y(_17321_));
 sky130_fd_sc_hd__o211ai_2 _27205_ (.A1(_17261_),
    .A2(_17110_),
    .B1(_17318_),
    .C1(_17321_),
    .Y(_17322_));
 sky130_fd_sc_hd__a211o_2 _27206_ (.A1(_17318_),
    .A2(_17321_),
    .B1(_17261_),
    .C1(_17110_),
    .X(_17323_));
 sky130_fd_sc_hd__inv_2 _27207_ (.A(_17138_),
    .Y(_17324_));
 sky130_fd_sc_hd__and4_2 _27208_ (.A(iX[34]),
    .B(iX[35]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_17325_));
 sky130_fd_sc_hd__a22oi_2 _27209_ (.A1(iX[35]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[34]),
    .Y(_17326_));
 sky130_fd_sc_hd__nor2_2 _27210_ (.A(_17325_),
    .B(_17326_),
    .Y(_17327_));
 sky130_fd_sc_hd__nand2_2 _27211_ (.A(iX[33]),
    .B(iY[52]),
    .Y(_17328_));
 sky130_fd_sc_hd__xnor2_2 _27212_ (.A(_17327_),
    .B(_17328_),
    .Y(_17329_));
 sky130_fd_sc_hd__o21ba_2 _27213_ (.A1(_17116_),
    .A2(_17118_),
    .B1_N(_17115_),
    .X(_17331_));
 sky130_fd_sc_hd__xnor2_2 _27214_ (.A(_17329_),
    .B(_17331_),
    .Y(_17332_));
 sky130_fd_sc_hd__nand2_2 _27215_ (.A(iX[32]),
    .B(iY[53]),
    .Y(_17333_));
 sky130_fd_sc_hd__xor2_2 _27216_ (.A(_17332_),
    .B(_17333_),
    .X(_17334_));
 sky130_fd_sc_hd__or3_2 _27217_ (.A(_17126_),
    .B(_17130_),
    .C(_17131_),
    .X(_17335_));
 sky130_fd_sc_hd__o21ba_2 _27218_ (.A1(_17055_),
    .A2(_17058_),
    .B1_N(_17054_),
    .X(_17336_));
 sky130_fd_sc_hd__and4_2 _27219_ (.A(iX[37]),
    .B(iX[38]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_17337_));
 sky130_fd_sc_hd__a22oi_2 _27220_ (.A1(iX[38]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[37]),
    .Y(_17338_));
 sky130_fd_sc_hd__nor2_2 _27221_ (.A(_17337_),
    .B(_17338_),
    .Y(_17339_));
 sky130_fd_sc_hd__nand2_2 _27222_ (.A(iX[36]),
    .B(iY[49]),
    .Y(_17340_));
 sky130_fd_sc_hd__xnor2_2 _27223_ (.A(_17339_),
    .B(_17340_),
    .Y(_17342_));
 sky130_fd_sc_hd__xnor2_2 _27224_ (.A(_17336_),
    .B(_17342_),
    .Y(_17343_));
 sky130_fd_sc_hd__o21ai_2 _27225_ (.A1(_17127_),
    .A2(_17131_),
    .B1(_17343_),
    .Y(_17344_));
 sky130_fd_sc_hd__or3_2 _27226_ (.A(_17127_),
    .B(_17131_),
    .C(_17343_),
    .X(_17345_));
 sky130_fd_sc_hd__nand2_2 _27227_ (.A(_17344_),
    .B(_17345_),
    .Y(_17346_));
 sky130_fd_sc_hd__a21oi_2 _27228_ (.A1(_17335_),
    .A2(_17135_),
    .B1(_17346_),
    .Y(_17347_));
 sky130_fd_sc_hd__and3_2 _27229_ (.A(_17335_),
    .B(_17135_),
    .C(_17346_),
    .X(_17348_));
 sky130_fd_sc_hd__or3_2 _27230_ (.A(_17334_),
    .B(_17347_),
    .C(_17348_),
    .X(_17349_));
 sky130_fd_sc_hd__o21ai_2 _27231_ (.A1(_17347_),
    .A2(_17348_),
    .B1(_17334_),
    .Y(_17350_));
 sky130_fd_sc_hd__nand2_2 _27232_ (.A(_17349_),
    .B(_17350_),
    .Y(_17351_));
 sky130_fd_sc_hd__a21oi_2 _27233_ (.A1(_17071_),
    .A2(_17073_),
    .B1(_17351_),
    .Y(_17353_));
 sky130_fd_sc_hd__and3_2 _27234_ (.A(_17071_),
    .B(_17073_),
    .C(_17351_),
    .X(_17354_));
 sky130_fd_sc_hd__a211oi_2 _27235_ (.A1(_17324_),
    .A2(_17140_),
    .B1(_17353_),
    .C1(_17354_),
    .Y(_17355_));
 sky130_fd_sc_hd__o211a_2 _27236_ (.A1(_17353_),
    .A2(_17354_),
    .B1(_17324_),
    .C1(_17140_),
    .X(_17356_));
 sky130_fd_sc_hd__nor2_2 _27237_ (.A(_17355_),
    .B(_17356_),
    .Y(_17357_));
 sky130_fd_sc_hd__nand3_2 _27238_ (.A(_17322_),
    .B(_17323_),
    .C(_17357_),
    .Y(_17358_));
 sky130_fd_sc_hd__a21o_2 _27239_ (.A1(_17322_),
    .A2(_17323_),
    .B1(_17357_),
    .X(_17359_));
 sky130_fd_sc_hd__o211ai_2 _27240_ (.A1(_17113_),
    .A2(_17148_),
    .B1(_17358_),
    .C1(_17359_),
    .Y(_17360_));
 sky130_fd_sc_hd__a211o_2 _27241_ (.A1(_17358_),
    .A2(_17359_),
    .B1(_17113_),
    .C1(_17148_),
    .X(_17361_));
 sky130_fd_sc_hd__o21ai_2 _27242_ (.A1(_17143_),
    .A2(_17146_),
    .B1(_17120_),
    .Y(_17362_));
 sky130_fd_sc_hd__or3_2 _27243_ (.A(_17120_),
    .B(_17143_),
    .C(_17146_),
    .X(_17364_));
 sky130_fd_sc_hd__and2_2 _27244_ (.A(_17362_),
    .B(_17364_),
    .X(_17365_));
 sky130_fd_sc_hd__and3_2 _27245_ (.A(_17360_),
    .B(_17361_),
    .C(_17365_),
    .X(_17366_));
 sky130_fd_sc_hd__a21oi_2 _27246_ (.A1(_17360_),
    .A2(_17361_),
    .B1(_17365_),
    .Y(_17367_));
 sky130_fd_sc_hd__or2_2 _27247_ (.A(_17366_),
    .B(_17367_),
    .X(_17368_));
 sky130_fd_sc_hd__o21ba_2 _27248_ (.A1(_17151_),
    .A2(_17152_),
    .B1_N(_17150_),
    .X(_17369_));
 sky130_fd_sc_hd__xnor2_2 _27249_ (.A(_17368_),
    .B(_17369_),
    .Y(_17370_));
 sky130_fd_sc_hd__xnor2_2 _27250_ (.A(_17157_),
    .B(_17370_),
    .Y(_17371_));
 sky130_fd_sc_hd__xnor2_2 _27251_ (.A(_17159_),
    .B(_17371_),
    .Y(_17372_));
 sky130_fd_sc_hd__nor3_2 _27252_ (.A(_17260_),
    .B(_17169_),
    .C(_17372_),
    .Y(_17373_));
 sky130_fd_sc_hd__o21a_2 _27253_ (.A1(_17260_),
    .A2(_17169_),
    .B1(_17372_),
    .X(_17375_));
 sky130_fd_sc_hd__nor2_2 _27254_ (.A(_17373_),
    .B(_17375_),
    .Y(_17376_));
 sky130_fd_sc_hd__and2_2 _27255_ (.A(_16901_),
    .B(_17042_),
    .X(_17377_));
 sky130_fd_sc_hd__or2_2 _27256_ (.A(_17039_),
    .B(_17041_),
    .X(_17378_));
 sky130_fd_sc_hd__or2b_2 _27257_ (.A(_16949_),
    .B_N(_16906_),
    .X(_17379_));
 sky130_fd_sc_hd__o21a_2 _27258_ (.A1(_16905_),
    .A2(_16950_),
    .B1(_17379_),
    .X(_17380_));
 sky130_fd_sc_hd__xnor2_2 _27259_ (.A(_16928_),
    .B(_17380_),
    .Y(_17381_));
 sky130_fd_sc_hd__nor2_2 _27260_ (.A(_17027_),
    .B(_17029_),
    .Y(_17382_));
 sky130_fd_sc_hd__and2_2 _27261_ (.A(_16951_),
    .B(_17030_),
    .X(_17383_));
 sky130_fd_sc_hd__or2_2 _27262_ (.A(_16944_),
    .B(_16946_),
    .X(_17384_));
 sky130_fd_sc_hd__nand2_2 _27263_ (.A(_16930_),
    .B(_16948_),
    .Y(_17386_));
 sky130_fd_sc_hd__nand2_2 _27264_ (.A(_16955_),
    .B(_16967_),
    .Y(_17387_));
 sky130_fd_sc_hd__nand2b_2 _27265_ (.A_N(_16969_),
    .B(_16953_),
    .Y(_17388_));
 sky130_fd_sc_hd__and3_2 _27266_ (.A(_14388_),
    .B(_16612_),
    .C(_16907_),
    .X(_17389_));
 sky130_fd_sc_hd__o22a_2 _27267_ (.A1(_15167_),
    .A2(_16255_),
    .B1(_16616_),
    .B2(_12468_),
    .X(_17390_));
 sky130_fd_sc_hd__or4_2 _27268_ (.A(_11570_),
    .B(_16922_),
    .C(_17389_),
    .D(_17390_),
    .X(_17391_));
 sky130_fd_sc_hd__buf_1 _27269_ (.A(_12838_),
    .X(_17392_));
 sky130_fd_sc_hd__inv_2 _27270_ (.A(_16921_),
    .Y(_17393_));
 sky130_fd_sc_hd__buf_1 _27271_ (.A(_17393_),
    .X(_17394_));
 sky130_fd_sc_hd__a2bb2o_2 _27272_ (.A1_N(_17389_),
    .A2_N(_17390_),
    .B1(_17392_),
    .B2(_17394_),
    .X(_17395_));
 sky130_fd_sc_hd__a21bo_2 _27273_ (.A1(_16909_),
    .A2(_16923_),
    .B1_N(_16908_),
    .X(_17397_));
 sky130_fd_sc_hd__nand3_2 _27274_ (.A(_17391_),
    .B(_17395_),
    .C(_17397_),
    .Y(_17398_));
 sky130_fd_sc_hd__a21o_2 _27275_ (.A1(_17391_),
    .A2(_17395_),
    .B1(_17397_),
    .X(_17399_));
 sky130_fd_sc_hd__a21o_2 _27276_ (.A1(_16912_),
    .A2(_16916_),
    .B1(_16920_),
    .X(_17400_));
 sky130_fd_sc_hd__nor2_2 _27277_ (.A(iY[21]),
    .B(iY[53]),
    .Y(_17401_));
 sky130_fd_sc_hd__nand2_2 _27278_ (.A(iY[21]),
    .B(iY[53]),
    .Y(_17402_));
 sky130_fd_sc_hd__or2b_2 _27279_ (.A(_17401_),
    .B_N(_17402_),
    .X(_17403_));
 sky130_fd_sc_hd__and3_4 _27280_ (.A(_16918_),
    .B(_17400_),
    .C(_17403_),
    .X(_17404_));
 sky130_fd_sc_hd__a21oi_2 _27281_ (.A1(_16918_),
    .A2(_17400_),
    .B1(_17403_),
    .Y(_17405_));
 sky130_fd_sc_hd__or2_2 _27282_ (.A(_17404_),
    .B(_17405_),
    .X(_17406_));
 sky130_fd_sc_hd__buf_6 _27283_ (.A(_17406_),
    .X(_17408_));
 sky130_fd_sc_hd__buf_6 _27284_ (.A(_17408_),
    .X(_17409_));
 sky130_fd_sc_hd__nor2_2 _27285_ (.A(_11579_),
    .B(_17409_),
    .Y(_17410_));
 sky130_fd_sc_hd__and3_2 _27286_ (.A(_17398_),
    .B(_17399_),
    .C(_17410_),
    .X(_17411_));
 sky130_fd_sc_hd__a21oi_2 _27287_ (.A1(_17398_),
    .A2(_17399_),
    .B1(_17410_),
    .Y(_17412_));
 sky130_fd_sc_hd__nand2_2 _27288_ (.A(_16935_),
    .B(_16938_),
    .Y(_17413_));
 sky130_fd_sc_hd__a21o_2 _27289_ (.A1(_16957_),
    .A2(_16959_),
    .B1(_16956_),
    .X(_17414_));
 sky130_fd_sc_hd__nor2_2 _27290_ (.A(_14343_),
    .B(_15596_),
    .Y(_17415_));
 sky130_fd_sc_hd__or3b_2 _27291_ (.A(_14640_),
    .B(_16237_),
    .C_N(_17415_),
    .X(_17416_));
 sky130_fd_sc_hd__a2bb2o_2 _27292_ (.A1_N(_14640_),
    .A2_N(_15597_),
    .B1(_15585_),
    .B2(_12816_),
    .X(_17417_));
 sky130_fd_sc_hd__nand4_2 _27293_ (.A(_14628_),
    .B(_16934_),
    .C(_17416_),
    .D(_17417_),
    .Y(_17419_));
 sky130_fd_sc_hd__a22o_2 _27294_ (.A1(_14628_),
    .A2(_16933_),
    .B1(_17416_),
    .B2(_17417_),
    .X(_17420_));
 sky130_fd_sc_hd__nand3_2 _27295_ (.A(_17414_),
    .B(_17419_),
    .C(_17420_),
    .Y(_17421_));
 sky130_fd_sc_hd__a21o_2 _27296_ (.A1(_17419_),
    .A2(_17420_),
    .B1(_17414_),
    .X(_17422_));
 sky130_fd_sc_hd__nand3_2 _27297_ (.A(_17413_),
    .B(_17421_),
    .C(_17422_),
    .Y(_17423_));
 sky130_fd_sc_hd__a21o_2 _27298_ (.A1(_17421_),
    .A2(_17422_),
    .B1(_17413_),
    .X(_17424_));
 sky130_fd_sc_hd__a21bo_2 _27299_ (.A1(_16931_),
    .A2(_16941_),
    .B1_N(_16940_),
    .X(_17425_));
 sky130_fd_sc_hd__and3_2 _27300_ (.A(_17423_),
    .B(_17424_),
    .C(_17425_),
    .X(_17426_));
 sky130_fd_sc_hd__a21oi_2 _27301_ (.A1(_17423_),
    .A2(_17424_),
    .B1(_17425_),
    .Y(_17427_));
 sky130_fd_sc_hd__nor4_2 _27302_ (.A(_17411_),
    .B(_17412_),
    .C(_17426_),
    .D(_17427_),
    .Y(_17428_));
 sky130_fd_sc_hd__o22a_2 _27303_ (.A1(_17411_),
    .A2(_17412_),
    .B1(_17426_),
    .B2(_17427_),
    .X(_17430_));
 sky130_fd_sc_hd__a211oi_2 _27304_ (.A1(_17387_),
    .A2(_17388_),
    .B1(_17428_),
    .C1(_17430_),
    .Y(_17431_));
 sky130_fd_sc_hd__o211a_2 _27305_ (.A1(_17428_),
    .A2(_17430_),
    .B1(_17387_),
    .C1(_17388_),
    .X(_17432_));
 sky130_fd_sc_hd__a211oi_2 _27306_ (.A1(_17384_),
    .A2(_17386_),
    .B1(_17431_),
    .C1(_17432_),
    .Y(_17433_));
 sky130_fd_sc_hd__o211a_2 _27307_ (.A1(_17431_),
    .A2(_17432_),
    .B1(_17384_),
    .C1(_17386_),
    .X(_17434_));
 sky130_fd_sc_hd__nor2_2 _27308_ (.A(_17433_),
    .B(_17434_),
    .Y(_17435_));
 sky130_fd_sc_hd__or2_2 _27309_ (.A(_16964_),
    .B(_16965_),
    .X(_17436_));
 sky130_fd_sc_hd__o21ai_2 _27310_ (.A1(_16960_),
    .A2(_16966_),
    .B1(_17436_),
    .Y(_17437_));
 sky130_fd_sc_hd__and2b_2 _27311_ (.A_N(_16978_),
    .B(_16973_),
    .X(_17438_));
 sky130_fd_sc_hd__a21o_2 _27312_ (.A1(_16972_),
    .A2(_16980_),
    .B1(_17438_),
    .X(_17439_));
 sky130_fd_sc_hd__nand2_2 _27313_ (.A(_14652_),
    .B(_14605_),
    .Y(_17441_));
 sky130_fd_sc_hd__nand2_2 _27314_ (.A(_14648_),
    .B(_14410_),
    .Y(_17442_));
 sky130_fd_sc_hd__xor2_2 _27315_ (.A(_17441_),
    .B(_17442_),
    .X(_17443_));
 sky130_fd_sc_hd__nor2_2 _27316_ (.A(_14357_),
    .B(_15173_),
    .Y(_17444_));
 sky130_fd_sc_hd__xnor2_2 _27317_ (.A(_17443_),
    .B(_17444_),
    .Y(_17445_));
 sky130_fd_sc_hd__nor2_2 _27318_ (.A(_13893_),
    .B(_14987_),
    .Y(_17446_));
 sky130_fd_sc_hd__o22a_2 _27319_ (.A1(_13891_),
    .A2(_13934_),
    .B1(_14987_),
    .B2(_14386_),
    .X(_17447_));
 sky130_fd_sc_hd__a31o_2 _27320_ (.A1(_13543_),
    .A2(_13938_),
    .A3(_17446_),
    .B1(_17447_),
    .X(_17448_));
 sky130_fd_sc_hd__nand2_2 _27321_ (.A(_13845_),
    .B(_14392_),
    .Y(_17449_));
 sky130_fd_sc_hd__xnor2_2 _27322_ (.A(_17448_),
    .B(_17449_),
    .Y(_17450_));
 sky130_fd_sc_hd__o22a_2 _27323_ (.A1(_16647_),
    .A2(_16961_),
    .B1(_16962_),
    .B2(_16963_),
    .X(_17452_));
 sky130_fd_sc_hd__xnor2_2 _27324_ (.A(_17450_),
    .B(_17452_),
    .Y(_17453_));
 sky130_fd_sc_hd__xor2_2 _27325_ (.A(_17445_),
    .B(_17453_),
    .X(_17454_));
 sky130_fd_sc_hd__xor2_2 _27326_ (.A(_17439_),
    .B(_17454_),
    .X(_17455_));
 sky130_fd_sc_hd__xnor2_2 _27327_ (.A(_17437_),
    .B(_17455_),
    .Y(_17456_));
 sky130_fd_sc_hd__nor3_2 _27328_ (.A(_16981_),
    .B(_17018_),
    .C(_17019_),
    .Y(_17457_));
 sky130_fd_sc_hd__and2_2 _27329_ (.A(_16976_),
    .B(_16977_),
    .X(_17458_));
 sky130_fd_sc_hd__a31o_2 _27330_ (.A1(_14637_),
    .A2(_16292_),
    .A3(_16975_),
    .B1(_17458_),
    .X(_17459_));
 sky130_fd_sc_hd__nor2_2 _27331_ (.A(_15219_),
    .B(_15220_),
    .Y(_17460_));
 sky130_fd_sc_hd__a31o_2 _27332_ (.A1(_12759_),
    .A2(_17460_),
    .A3(_16984_),
    .B1(_16982_),
    .X(_17461_));
 sky130_fd_sc_hd__buf_1 _27333_ (.A(_13274_),
    .X(_17463_));
 sky130_fd_sc_hd__or4b_2 _27334_ (.A(_12850_),
    .B(_15219_),
    .C(_15220_),
    .D_N(_16975_),
    .X(_17464_));
 sky130_fd_sc_hd__a32o_2 _27335_ (.A1(_14634_),
    .A2(_15223_),
    .A3(_15225_),
    .B1(_12846_),
    .B2(_15679_),
    .X(_17465_));
 sky130_fd_sc_hd__nand4_2 _27336_ (.A(_17463_),
    .B(_16292_),
    .C(_17464_),
    .D(_17465_),
    .Y(_17466_));
 sky130_fd_sc_hd__a22o_2 _27337_ (.A1(_17463_),
    .A2(_16292_),
    .B1(_17464_),
    .B2(_17465_),
    .X(_17467_));
 sky130_fd_sc_hd__nand3_2 _27338_ (.A(_17461_),
    .B(_17466_),
    .C(_17467_),
    .Y(_17468_));
 sky130_fd_sc_hd__a21o_2 _27339_ (.A1(_17466_),
    .A2(_17467_),
    .B1(_17461_),
    .X(_17469_));
 sky130_fd_sc_hd__and3_2 _27340_ (.A(_17459_),
    .B(_17468_),
    .C(_17469_),
    .X(_17470_));
 sky130_fd_sc_hd__a21oi_2 _27341_ (.A1(_17468_),
    .A2(_17469_),
    .B1(_17459_),
    .Y(_17471_));
 sky130_fd_sc_hd__or3b_2 _27342_ (.A(_12248_),
    .B(_16988_),
    .C_N(_16983_),
    .X(_17472_));
 sky130_fd_sc_hd__a22o_2 _27343_ (.A1(_12242_),
    .A2(_15900_),
    .B1(_16682_),
    .B2(_11842_),
    .X(_17474_));
 sky130_fd_sc_hd__nand2_2 _27344_ (.A(_17472_),
    .B(_17474_),
    .Y(_17475_));
 sky130_fd_sc_hd__nor2_2 _27345_ (.A(_14356_),
    .B(_16312_),
    .Y(_17476_));
 sky130_fd_sc_hd__xnor2_2 _27346_ (.A(_17475_),
    .B(_17476_),
    .Y(_17477_));
 sky130_fd_sc_hd__nand2_2 _27347_ (.A(iX[21]),
    .B(iX[53]),
    .Y(_17478_));
 sky130_fd_sc_hd__or2_2 _27348_ (.A(iX[21]),
    .B(iX[53]),
    .X(_17479_));
 sky130_fd_sc_hd__nand2_2 _27349_ (.A(_17478_),
    .B(_17479_),
    .Y(_17480_));
 sky130_fd_sc_hd__o21ba_2 _27350_ (.A1(_16993_),
    .A2(_16998_),
    .B1_N(_16989_),
    .X(_17481_));
 sky130_fd_sc_hd__xnor2_2 _27351_ (.A(_17480_),
    .B(_17481_),
    .Y(_17482_));
 sky130_fd_sc_hd__or4_4 _27352_ (.A(_11565_),
    .B(_11575_),
    .C(_16999_),
    .D(_17482_),
    .X(_17483_));
 sky130_fd_sc_hd__xor2_2 _27353_ (.A(_17480_),
    .B(_17481_),
    .X(_17485_));
 sky130_fd_sc_hd__a21o_2 _27354_ (.A1(_11381_),
    .A2(_17485_),
    .B1(_17000_),
    .X(_17486_));
 sky130_fd_sc_hd__nand4_2 _27355_ (.A(_15675_),
    .B(_16680_),
    .C(_17483_),
    .D(_17486_),
    .Y(_17487_));
 sky130_fd_sc_hd__buf_2 _27356_ (.A(_16680_),
    .X(_17488_));
 sky130_fd_sc_hd__a22o_2 _27357_ (.A1(_15675_),
    .A2(_17488_),
    .B1(_17483_),
    .B2(_17486_),
    .X(_17489_));
 sky130_fd_sc_hd__a31o_2 _27358_ (.A1(_15675_),
    .A2(_17006_),
    .A3(_17004_),
    .B1(_17002_),
    .X(_17490_));
 sky130_fd_sc_hd__nand3_2 _27359_ (.A(_17487_),
    .B(_17489_),
    .C(_17490_),
    .Y(_17491_));
 sky130_fd_sc_hd__a21o_2 _27360_ (.A1(_17487_),
    .A2(_17489_),
    .B1(_17490_),
    .X(_17492_));
 sky130_fd_sc_hd__nand3_2 _27361_ (.A(_17477_),
    .B(_17491_),
    .C(_17492_),
    .Y(_17493_));
 sky130_fd_sc_hd__a21o_2 _27362_ (.A1(_17491_),
    .A2(_17492_),
    .B1(_17477_),
    .X(_17494_));
 sky130_fd_sc_hd__a21bo_2 _27363_ (.A1(_16987_),
    .A2(_17013_),
    .B1_N(_17011_),
    .X(_17496_));
 sky130_fd_sc_hd__nand3_2 _27364_ (.A(_17493_),
    .B(_17494_),
    .C(_17496_),
    .Y(_17497_));
 sky130_fd_sc_hd__a21o_2 _27365_ (.A1(_17493_),
    .A2(_17494_),
    .B1(_17496_),
    .X(_17498_));
 sky130_fd_sc_hd__nand4bb_2 _27366_ (.A_N(_17470_),
    .B_N(_17471_),
    .C(_17497_),
    .D(_17498_),
    .Y(_17499_));
 sky130_fd_sc_hd__a2bb2o_2 _27367_ (.A1_N(_17470_),
    .A2_N(_17471_),
    .B1(_17497_),
    .B2(_17498_),
    .X(_17500_));
 sky130_fd_sc_hd__o211a_2 _27368_ (.A1(_17018_),
    .A2(_17457_),
    .B1(_17499_),
    .C1(_17500_),
    .X(_17501_));
 sky130_fd_sc_hd__a211oi_2 _27369_ (.A1(_17499_),
    .A2(_17500_),
    .B1(_17018_),
    .C1(_17457_),
    .Y(_17502_));
 sky130_fd_sc_hd__nor3_2 _27370_ (.A(_17456_),
    .B(_17501_),
    .C(_17502_),
    .Y(_17503_));
 sky130_fd_sc_hd__o21a_2 _27371_ (.A1(_17501_),
    .A2(_17502_),
    .B1(_17456_),
    .X(_17504_));
 sky130_fd_sc_hd__o21ba_2 _27372_ (.A1(_16970_),
    .A2(_17024_),
    .B1_N(_17022_),
    .X(_17505_));
 sky130_fd_sc_hd__or3_4 _27373_ (.A(_17503_),
    .B(_17504_),
    .C(_17505_),
    .X(_17507_));
 sky130_fd_sc_hd__o21ai_2 _27374_ (.A1(_17503_),
    .A2(_17504_),
    .B1(_17505_),
    .Y(_17508_));
 sky130_fd_sc_hd__and2_4 _27375_ (.A(_17507_),
    .B(_17508_),
    .X(_17509_));
 sky130_fd_sc_hd__xnor2_2 _27376_ (.A(_17435_),
    .B(_17509_),
    .Y(_17510_));
 sky130_fd_sc_hd__o21ba_2 _27377_ (.A1(_17382_),
    .A2(_17383_),
    .B1_N(_17510_),
    .X(_17511_));
 sky130_fd_sc_hd__or3b_2 _27378_ (.A(_17382_),
    .B(_17383_),
    .C_N(_17510_),
    .X(_17512_));
 sky130_fd_sc_hd__nand2b_2 _27379_ (.A_N(_17511_),
    .B(_17512_),
    .Y(_17513_));
 sky130_fd_sc_hd__xor2_2 _27380_ (.A(_17381_),
    .B(_17513_),
    .X(_17514_));
 sky130_fd_sc_hd__a21o_2 _27381_ (.A1(_16904_),
    .A2(_17037_),
    .B1(_17036_),
    .X(_17515_));
 sky130_fd_sc_hd__xor2_2 _27382_ (.A(_17514_),
    .B(_17515_),
    .X(_17516_));
 sky130_fd_sc_hd__xor2_2 _27383_ (.A(_17378_),
    .B(_17516_),
    .X(_17518_));
 sky130_fd_sc_hd__xnor2_2 _27384_ (.A(_17377_),
    .B(_17518_),
    .Y(_17519_));
 sky130_fd_sc_hd__inv_2 _27385_ (.A(_17519_),
    .Y(_17520_));
 sky130_fd_sc_hd__a31oi_2 _27386_ (.A1(_15579_),
    .A2(_16893_),
    .A3(_16894_),
    .B1(_16899_),
    .Y(_17521_));
 sky130_fd_sc_hd__inv_2 _27387_ (.A(_17044_),
    .Y(_17522_));
 sky130_fd_sc_hd__or2b_2 _27388_ (.A(_16895_),
    .B_N(_17043_),
    .X(_17523_));
 sky130_fd_sc_hd__o21a_2 _27389_ (.A1(_17521_),
    .A2(_17522_),
    .B1(_17523_),
    .X(_17524_));
 sky130_fd_sc_hd__xnor2_2 _27390_ (.A(_17520_),
    .B(_17524_),
    .Y(_17525_));
 sky130_fd_sc_hd__xnor2_2 _27391_ (.A(_17376_),
    .B(_17525_),
    .Y(_17526_));
 sky130_fd_sc_hd__xnor2_2 _27392_ (.A(oO[21]),
    .B(_17526_),
    .Y(_17527_));
 sky130_fd_sc_hd__o21a_2 _27393_ (.A1(oO[20]),
    .A2(_17174_),
    .B1(_17173_),
    .X(_17529_));
 sky130_fd_sc_hd__xnor2_2 _27394_ (.A(_17527_),
    .B(_17529_),
    .Y(_17530_));
 sky130_fd_sc_hd__nor2_2 _27395_ (.A(_17175_),
    .B(_17179_),
    .Y(_17531_));
 sky130_fd_sc_hd__nor2_2 _27396_ (.A(_17531_),
    .B(_17181_),
    .Y(_17532_));
 sky130_fd_sc_hd__xor2_2 _27397_ (.A(_17530_),
    .B(_17532_),
    .X(_17533_));
 sky130_fd_sc_hd__and2_2 _27398_ (.A(_17259_),
    .B(_17533_),
    .X(_17534_));
 sky130_fd_sc_hd__nor2_2 _27399_ (.A(_17259_),
    .B(_17533_),
    .Y(_17535_));
 sky130_fd_sc_hd__nor2_2 _27400_ (.A(_17534_),
    .B(_17535_),
    .Y(_17536_));
 sky130_fd_sc_hd__and2b_2 _27401_ (.A_N(_16890_),
    .B(_17183_),
    .X(_17537_));
 sky130_fd_sc_hd__and2b_2 _27402_ (.A_N(_17184_),
    .B(_17190_),
    .X(_17538_));
 sky130_fd_sc_hd__nor2_2 _27403_ (.A(_17537_),
    .B(_17538_),
    .Y(_17540_));
 sky130_fd_sc_hd__xnor2_2 _27404_ (.A(_17536_),
    .B(_17540_),
    .Y(oO[53]));
 sky130_fd_sc_hd__o21ai_2 _27405_ (.A1(_16844_),
    .A2(_16865_),
    .B1(_17241_),
    .Y(_17541_));
 sky130_fd_sc_hd__nand2_2 _27406_ (.A(iY[23]),
    .B(iX[31]),
    .Y(_17542_));
 sky130_fd_sc_hd__and2_2 _27407_ (.A(iY[25]),
    .B(iX[30]),
    .X(_17543_));
 sky130_fd_sc_hd__and3_2 _27408_ (.A(iY[24]),
    .B(iX[29]),
    .C(_17543_),
    .X(_17544_));
 sky130_fd_sc_hd__a22oi_2 _27409_ (.A1(iY[25]),
    .A2(iX[29]),
    .B1(iX[30]),
    .B2(iY[24]),
    .Y(_17545_));
 sky130_fd_sc_hd__and4bb_2 _27410_ (.A_N(_17544_),
    .B_N(_17545_),
    .C(iY[26]),
    .D(iX[28]),
    .X(_17546_));
 sky130_fd_sc_hd__o2bb2a_2 _27411_ (.A1_N(iY[26]),
    .A2_N(iX[28]),
    .B1(_17544_),
    .B2(_17545_),
    .X(_17547_));
 sky130_fd_sc_hd__nor2_2 _27412_ (.A(_17546_),
    .B(_17547_),
    .Y(_17548_));
 sky130_fd_sc_hd__xnor2_2 _27413_ (.A(_17195_),
    .B(_17548_),
    .Y(_17550_));
 sky130_fd_sc_hd__a31o_2 _27414_ (.A1(iY[26]),
    .A2(iX[27]),
    .A3(_17202_),
    .B1(_17200_),
    .X(_17551_));
 sky130_fd_sc_hd__and2b_2 _27415_ (.A_N(_17550_),
    .B(_17551_),
    .X(_17552_));
 sky130_fd_sc_hd__and2b_2 _27416_ (.A_N(_17551_),
    .B(_17550_),
    .X(_17553_));
 sky130_fd_sc_hd__or2_2 _27417_ (.A(_17552_),
    .B(_17553_),
    .X(_17554_));
 sky130_fd_sc_hd__a21oi_2 _27418_ (.A1(_17205_),
    .A2(_17208_),
    .B1(_17554_),
    .Y(_17555_));
 sky130_fd_sc_hd__and3_2 _27419_ (.A(_17205_),
    .B(_17208_),
    .C(_17554_),
    .X(_17556_));
 sky130_fd_sc_hd__or3_2 _27420_ (.A(_17213_),
    .B(_17555_),
    .C(_17556_),
    .X(_17557_));
 sky130_fd_sc_hd__o21ai_2 _27421_ (.A1(_17555_),
    .A2(_17556_),
    .B1(_17213_),
    .Y(_17558_));
 sky130_fd_sc_hd__or2b_2 _27422_ (.A(_17228_),
    .B_N(_17227_),
    .X(_17559_));
 sky130_fd_sc_hd__and4_2 _27423_ (.A(iX[26]),
    .B(iX[27]),
    .C(iY[27]),
    .D(iY[28]),
    .X(_17561_));
 sky130_fd_sc_hd__a22oi_2 _27424_ (.A1(iX[27]),
    .A2(iY[27]),
    .B1(iY[28]),
    .B2(iX[26]),
    .Y(_17562_));
 sky130_fd_sc_hd__nor2_2 _27425_ (.A(_17561_),
    .B(_17562_),
    .Y(_17563_));
 sky130_fd_sc_hd__nand2_2 _27426_ (.A(iX[25]),
    .B(iY[29]),
    .Y(_17564_));
 sky130_fd_sc_hd__xnor2_2 _27427_ (.A(_17563_),
    .B(_17564_),
    .Y(_17565_));
 sky130_fd_sc_hd__o21ba_2 _27428_ (.A1(_17224_),
    .A2(_17226_),
    .B1_N(_17223_),
    .X(_17566_));
 sky130_fd_sc_hd__xnor2_2 _27429_ (.A(_17565_),
    .B(_17566_),
    .Y(_17567_));
 sky130_fd_sc_hd__nand3_2 _27430_ (.A(iX[24]),
    .B(iY[30]),
    .C(_17567_),
    .Y(_17568_));
 sky130_fd_sc_hd__a21o_2 _27431_ (.A1(iX[24]),
    .A2(iY[30]),
    .B1(_17567_),
    .X(_17569_));
 sky130_fd_sc_hd__nand2_2 _27432_ (.A(_17568_),
    .B(_17569_),
    .Y(_17570_));
 sky130_fd_sc_hd__a21oi_2 _27433_ (.A1(_17559_),
    .A2(_17230_),
    .B1(_17570_),
    .Y(_17572_));
 sky130_fd_sc_hd__and3_2 _27434_ (.A(_17559_),
    .B(_17230_),
    .C(_17570_),
    .X(_17573_));
 sky130_fd_sc_hd__nor2_2 _27435_ (.A(_17572_),
    .B(_17573_),
    .Y(_17574_));
 sky130_fd_sc_hd__nand2_2 _27436_ (.A(iX[23]),
    .B(iY[31]),
    .Y(_17575_));
 sky130_fd_sc_hd__xnor2_2 _27437_ (.A(_17574_),
    .B(_17575_),
    .Y(_17576_));
 sky130_fd_sc_hd__and3_2 _27438_ (.A(_17557_),
    .B(_17558_),
    .C(_17576_),
    .X(_17577_));
 sky130_fd_sc_hd__a21oi_2 _27439_ (.A1(_17557_),
    .A2(_17558_),
    .B1(_17576_),
    .Y(_17578_));
 sky130_fd_sc_hd__or2_2 _27440_ (.A(_17577_),
    .B(_17578_),
    .X(_17579_));
 sky130_fd_sc_hd__a21o_2 _27441_ (.A1(_17218_),
    .A2(_17239_),
    .B1(_17579_),
    .X(_17580_));
 sky130_fd_sc_hd__nand3_2 _27442_ (.A(_17218_),
    .B(_17239_),
    .C(_17579_),
    .Y(_17581_));
 sky130_fd_sc_hd__nand2_2 _27443_ (.A(_17580_),
    .B(_17581_),
    .Y(_17583_));
 sky130_fd_sc_hd__xor2_2 _27444_ (.A(_17542_),
    .B(_17583_),
    .X(_17584_));
 sky130_fd_sc_hd__nand2_2 _27445_ (.A(_17245_),
    .B(_17584_),
    .Y(_17585_));
 sky130_fd_sc_hd__or2_2 _27446_ (.A(_17245_),
    .B(_17584_),
    .X(_17586_));
 sky130_fd_sc_hd__nand2_2 _27447_ (.A(_17585_),
    .B(_17586_),
    .Y(_17587_));
 sky130_fd_sc_hd__xnor2_2 _27448_ (.A(_17541_),
    .B(_17587_),
    .Y(_17588_));
 sky130_fd_sc_hd__inv_2 _27449_ (.A(_16867_),
    .Y(_17589_));
 sky130_fd_sc_hd__o21ai_2 _27450_ (.A1(_17589_),
    .A2(_16871_),
    .B1(_17247_),
    .Y(_17590_));
 sky130_fd_sc_hd__or2_2 _27451_ (.A(_17588_),
    .B(_17590_),
    .X(_17591_));
 sky130_fd_sc_hd__nand2_2 _27452_ (.A(_17588_),
    .B(_17590_),
    .Y(_17592_));
 sky130_fd_sc_hd__nand2_2 _27453_ (.A(_17591_),
    .B(_17592_),
    .Y(_17594_));
 sky130_fd_sc_hd__o21ba_2 _27454_ (.A1(_17235_),
    .A2(_17237_),
    .B1_N(_17234_),
    .X(_17595_));
 sky130_fd_sc_hd__or2_2 _27455_ (.A(_17594_),
    .B(_17595_),
    .X(_17596_));
 sky130_fd_sc_hd__nand2_2 _27456_ (.A(_17594_),
    .B(_17595_),
    .Y(_17597_));
 sky130_fd_sc_hd__nand2_2 _27457_ (.A(_17596_),
    .B(_17597_),
    .Y(_17598_));
 sky130_fd_sc_hd__a21oi_2 _27458_ (.A1(_17251_),
    .A2(_17254_),
    .B1(_17250_),
    .Y(_17599_));
 sky130_fd_sc_hd__or2_2 _27459_ (.A(_17598_),
    .B(_17599_),
    .X(_17600_));
 sky130_fd_sc_hd__nand2_2 _27460_ (.A(_17598_),
    .B(_17599_),
    .Y(_17601_));
 sky130_fd_sc_hd__nand2_2 _27461_ (.A(_17600_),
    .B(_17601_),
    .Y(_17602_));
 sky130_fd_sc_hd__a21oi_2 _27462_ (.A1(_17192_),
    .A2(_17258_),
    .B1(_17256_),
    .Y(_17603_));
 sky130_fd_sc_hd__xnor2_2 _27463_ (.A(_17602_),
    .B(_17603_),
    .Y(_17605_));
 sky130_fd_sc_hd__or2b_2 _27464_ (.A(_17376_),
    .B_N(_17525_),
    .X(_17606_));
 sky130_fd_sc_hd__or2b_2 _27465_ (.A(oO[21]),
    .B_N(_17526_),
    .X(_17607_));
 sky130_fd_sc_hd__nor2_2 _27466_ (.A(_17378_),
    .B(_17516_),
    .Y(_17608_));
 sky130_fd_sc_hd__nor2b_2 _27467_ (.A(_17514_),
    .B_N(_17515_),
    .Y(_17609_));
 sky130_fd_sc_hd__or3_2 _27468_ (.A(_16620_),
    .B(_16927_),
    .C(_17380_),
    .X(_17610_));
 sky130_fd_sc_hd__inv_2 _27469_ (.A(_17398_),
    .Y(_17611_));
 sky130_fd_sc_hd__nor2_2 _27470_ (.A(_17611_),
    .B(_17411_),
    .Y(_17612_));
 sky130_fd_sc_hd__o21ba_2 _27471_ (.A1(_17431_),
    .A2(_17433_),
    .B1_N(_17612_),
    .X(_17613_));
 sky130_fd_sc_hd__or3b_2 _27472_ (.A(_17431_),
    .B(_17433_),
    .C_N(_17612_),
    .X(_17614_));
 sky130_fd_sc_hd__or2b_2 _27473_ (.A(_17613_),
    .B_N(_17614_),
    .X(_17616_));
 sky130_fd_sc_hd__or2_2 _27474_ (.A(_17426_),
    .B(_17428_),
    .X(_17617_));
 sky130_fd_sc_hd__and2_2 _27475_ (.A(_17439_),
    .B(_17454_),
    .X(_17618_));
 sky130_fd_sc_hd__a21o_2 _27476_ (.A1(_17437_),
    .A2(_17455_),
    .B1(_17618_),
    .X(_17619_));
 sky130_fd_sc_hd__nand2_2 _27477_ (.A(iY[22]),
    .B(iY[54]),
    .Y(_17620_));
 sky130_fd_sc_hd__or2_2 _27478_ (.A(iY[22]),
    .B(iY[54]),
    .X(_17621_));
 sky130_fd_sc_hd__nand2_2 _27479_ (.A(_17620_),
    .B(_17621_),
    .Y(_17622_));
 sky130_fd_sc_hd__a311oi_4 _27480_ (.A1(_16918_),
    .A2(_17400_),
    .A3(_17402_),
    .B1(_17622_),
    .C1(_17401_),
    .Y(_17623_));
 sky130_fd_sc_hd__a21o_2 _27481_ (.A1(_16918_),
    .A2(_17402_),
    .B1(_17401_),
    .X(_17624_));
 sky130_fd_sc_hd__o211a_2 _27482_ (.A1(_17400_),
    .A2(_17401_),
    .B1(_17622_),
    .C1(_17624_),
    .X(_17625_));
 sky130_fd_sc_hd__or2_4 _27483_ (.A(_17623_),
    .B(_17625_),
    .X(_17627_));
 sky130_fd_sc_hd__buf_2 _27484_ (.A(_17627_),
    .X(_17628_));
 sky130_fd_sc_hd__nor2_2 _27485_ (.A(_17404_),
    .B(_17405_),
    .Y(_17629_));
 sky130_fd_sc_hd__buf_6 _27486_ (.A(_17629_),
    .X(_17630_));
 sky130_fd_sc_hd__nand2_2 _27487_ (.A(_17392_),
    .B(_17630_),
    .Y(_17631_));
 sky130_fd_sc_hd__o21ai_2 _27488_ (.A1(_11579_),
    .A2(_17628_),
    .B1(_17631_),
    .Y(_17632_));
 sky130_fd_sc_hd__or3_2 _27489_ (.A(_11578_),
    .B(_17631_),
    .C(_17628_),
    .X(_17633_));
 sky130_fd_sc_hd__nand2_2 _27490_ (.A(_17632_),
    .B(_17633_),
    .Y(_17634_));
 sky130_fd_sc_hd__nor2_2 _27491_ (.A(_15167_),
    .B(_16617_),
    .Y(_17635_));
 sky130_fd_sc_hd__nor2_2 _27492_ (.A(_14346_),
    .B(_16257_),
    .Y(_17636_));
 sky130_fd_sc_hd__xnor2_2 _27493_ (.A(_17635_),
    .B(_17636_),
    .Y(_17638_));
 sky130_fd_sc_hd__or2_2 _27494_ (.A(_16625_),
    .B(_16922_),
    .X(_17639_));
 sky130_fd_sc_hd__xnor2_2 _27495_ (.A(_17638_),
    .B(_17639_),
    .Y(_17640_));
 sky130_fd_sc_hd__or2b_2 _27496_ (.A(_17389_),
    .B_N(_17391_),
    .X(_17641_));
 sky130_fd_sc_hd__xor2_2 _27497_ (.A(_17640_),
    .B(_17641_),
    .X(_17642_));
 sky130_fd_sc_hd__xnor2_2 _27498_ (.A(_17634_),
    .B(_17642_),
    .Y(_17643_));
 sky130_fd_sc_hd__nand2_2 _27499_ (.A(_17416_),
    .B(_17419_),
    .Y(_17644_));
 sky130_fd_sc_hd__nor2_2 _27500_ (.A(_17441_),
    .B(_17442_),
    .Y(_17645_));
 sky130_fd_sc_hd__a21o_2 _27501_ (.A1(_17443_),
    .A2(_17444_),
    .B1(_17645_),
    .X(_17646_));
 sky130_fd_sc_hd__or3b_2 _27502_ (.A(_14357_),
    .B(_16237_),
    .C_N(_17415_),
    .X(_17647_));
 sky130_fd_sc_hd__a21o_2 _27503_ (.A1(_16277_),
    .A2(_15585_),
    .B1(_17415_),
    .X(_17649_));
 sky130_fd_sc_hd__nand2_2 _27504_ (.A(_17647_),
    .B(_17649_),
    .Y(_17650_));
 sky130_fd_sc_hd__nor2_2 _27505_ (.A(_14640_),
    .B(_15834_),
    .Y(_17651_));
 sky130_fd_sc_hd__xnor2_2 _27506_ (.A(_17650_),
    .B(_17651_),
    .Y(_17652_));
 sky130_fd_sc_hd__xor2_2 _27507_ (.A(_17646_),
    .B(_17652_),
    .X(_17653_));
 sky130_fd_sc_hd__xnor2_2 _27508_ (.A(_17644_),
    .B(_17653_),
    .Y(_17654_));
 sky130_fd_sc_hd__and2_2 _27509_ (.A(_17421_),
    .B(_17423_),
    .X(_17655_));
 sky130_fd_sc_hd__xnor2_2 _27510_ (.A(_17654_),
    .B(_17655_),
    .Y(_17656_));
 sky130_fd_sc_hd__xor2_2 _27511_ (.A(_17643_),
    .B(_17656_),
    .X(_17657_));
 sky130_fd_sc_hd__xnor2_2 _27512_ (.A(_17619_),
    .B(_17657_),
    .Y(_17658_));
 sky130_fd_sc_hd__xnor2_2 _27513_ (.A(_17617_),
    .B(_17658_),
    .Y(_17660_));
 sky130_fd_sc_hd__or2_2 _27514_ (.A(_17445_),
    .B(_17453_),
    .X(_17661_));
 sky130_fd_sc_hd__o21ai_2 _27515_ (.A1(_17450_),
    .A2(_17452_),
    .B1(_17661_),
    .Y(_17662_));
 sky130_fd_sc_hd__and3_2 _27516_ (.A(_17461_),
    .B(_17466_),
    .C(_17467_),
    .X(_17663_));
 sky130_fd_sc_hd__nand2_2 _27517_ (.A(_13845_),
    .B(_14608_),
    .Y(_17664_));
 sky130_fd_sc_hd__a22o_2 _27518_ (.A1(_13845_),
    .A2(_14410_),
    .B1(_14605_),
    .B2(_14648_),
    .X(_17665_));
 sky130_fd_sc_hd__o21a_2 _27519_ (.A1(_17442_),
    .A2(_17664_),
    .B1(_17665_),
    .X(_17666_));
 sky130_fd_sc_hd__nor2_2 _27520_ (.A(_14352_),
    .B(_14948_),
    .Y(_17667_));
 sky130_fd_sc_hd__xnor2_2 _27521_ (.A(_17666_),
    .B(_17667_),
    .Y(_17668_));
 sky130_fd_sc_hd__nor2_2 _27522_ (.A(_14386_),
    .B(_15004_),
    .Y(_17669_));
 sky130_fd_sc_hd__xnor2_2 _27523_ (.A(_17446_),
    .B(_17669_),
    .Y(_17671_));
 sky130_fd_sc_hd__nand2_2 _27524_ (.A(_13938_),
    .B(_14391_),
    .Y(_17672_));
 sky130_fd_sc_hd__xnor2_2 _27525_ (.A(_17671_),
    .B(_17672_),
    .Y(_17673_));
 sky130_fd_sc_hd__nand2_2 _27526_ (.A(_13889_),
    .B(_15208_),
    .Y(_17674_));
 sky130_fd_sc_hd__o22a_2 _27527_ (.A1(_16961_),
    .A2(_17674_),
    .B1(_17447_),
    .B2(_17449_),
    .X(_17675_));
 sky130_fd_sc_hd__xnor2_2 _27528_ (.A(_17673_),
    .B(_17675_),
    .Y(_17676_));
 sky130_fd_sc_hd__xor2_2 _27529_ (.A(_17668_),
    .B(_17676_),
    .X(_17677_));
 sky130_fd_sc_hd__o21ai_2 _27530_ (.A1(_17663_),
    .A2(_17470_),
    .B1(_17677_),
    .Y(_17678_));
 sky130_fd_sc_hd__or3_4 _27531_ (.A(_17663_),
    .B(_17470_),
    .C(_17677_),
    .X(_17679_));
 sky130_fd_sc_hd__nand2_2 _27532_ (.A(_17678_),
    .B(_17679_),
    .Y(_17680_));
 sky130_fd_sc_hd__xnor2_2 _27533_ (.A(_17662_),
    .B(_17680_),
    .Y(_17682_));
 sky130_fd_sc_hd__nand2_2 _27534_ (.A(_17464_),
    .B(_17466_),
    .Y(_17683_));
 sky130_fd_sc_hd__a21bo_2 _27535_ (.A1(_17474_),
    .A2(_17476_),
    .B1_N(_17472_),
    .X(_17684_));
 sky130_fd_sc_hd__nor2_2 _27536_ (.A(_14641_),
    .B(_14998_),
    .Y(_17685_));
 sky130_fd_sc_hd__nor2_2 _27537_ (.A(_12849_),
    .B(_16312_),
    .Y(_17686_));
 sky130_fd_sc_hd__or4b_4 _27538_ (.A(_12773_),
    .B(_15219_),
    .C(_15220_),
    .D_N(_17686_),
    .X(_17687_));
 sky130_fd_sc_hd__a32o_2 _27539_ (.A1(_12846_),
    .A2(_15224_),
    .A3(_15226_),
    .B1(_15672_),
    .B2(_14634_),
    .X(_17688_));
 sky130_fd_sc_hd__nand3_2 _27540_ (.A(_17685_),
    .B(_17687_),
    .C(_17688_),
    .Y(_17689_));
 sky130_fd_sc_hd__a21o_2 _27541_ (.A1(_17687_),
    .A2(_17688_),
    .B1(_17685_),
    .X(_17690_));
 sky130_fd_sc_hd__and3_2 _27542_ (.A(_17684_),
    .B(_17689_),
    .C(_17690_),
    .X(_17691_));
 sky130_fd_sc_hd__a21o_2 _27543_ (.A1(_17689_),
    .A2(_17690_),
    .B1(_17684_),
    .X(_17693_));
 sky130_fd_sc_hd__nand2b_2 _27544_ (.A_N(_17691_),
    .B(_17693_),
    .Y(_17694_));
 sky130_fd_sc_hd__xnor2_2 _27545_ (.A(_17683_),
    .B(_17694_),
    .Y(_17695_));
 sky130_fd_sc_hd__buf_1 _27546_ (.A(_16677_),
    .X(_17696_));
 sky130_fd_sc_hd__nor2_2 _27547_ (.A(_15646_),
    .B(_17696_),
    .Y(_17697_));
 sky130_fd_sc_hd__nor2_2 _27548_ (.A(_15650_),
    .B(_16988_),
    .Y(_17698_));
 sky130_fd_sc_hd__o22a_2 _27549_ (.A1(_14978_),
    .A2(_16988_),
    .B1(_17007_),
    .B2(_15650_),
    .X(_17699_));
 sky130_fd_sc_hd__a31o_2 _27550_ (.A1(_14980_),
    .A2(_17488_),
    .A3(_17698_),
    .B1(_17699_),
    .X(_17700_));
 sky130_fd_sc_hd__xnor2_2 _27551_ (.A(_17697_),
    .B(_17700_),
    .Y(_17701_));
 sky130_fd_sc_hd__buf_1 _27552_ (.A(_17003_),
    .X(_17702_));
 sky130_fd_sc_hd__nand2_2 _27553_ (.A(_15675_),
    .B(_17702_),
    .Y(_17704_));
 sky130_fd_sc_hd__nand2_2 _27554_ (.A(_11585_),
    .B(_17485_),
    .Y(_17705_));
 sky130_fd_sc_hd__or2b_2 _27555_ (.A(_16989_),
    .B_N(_17478_),
    .X(_17706_));
 sky130_fd_sc_hd__o21bai_2 _27556_ (.A1(_16993_),
    .A2(_16998_),
    .B1_N(_17706_),
    .Y(_17707_));
 sky130_fd_sc_hd__and2_2 _27557_ (.A(iX[22]),
    .B(iX[54]),
    .X(_17708_));
 sky130_fd_sc_hd__nor2_2 _27558_ (.A(iX[22]),
    .B(iX[54]),
    .Y(_17709_));
 sky130_fd_sc_hd__nor2_2 _27559_ (.A(_17708_),
    .B(_17709_),
    .Y(_17710_));
 sky130_fd_sc_hd__and2_2 _27560_ (.A(_17479_),
    .B(_17710_),
    .X(_17711_));
 sky130_fd_sc_hd__nand2_2 _27561_ (.A(_17707_),
    .B(_17711_),
    .Y(_17712_));
 sky130_fd_sc_hd__a21o_2 _27562_ (.A1(_17479_),
    .A2(_17707_),
    .B1(_17710_),
    .X(_17713_));
 sky130_fd_sc_hd__and3_4 _27563_ (.A(_11380_),
    .B(_17712_),
    .C(_17713_),
    .X(_17715_));
 sky130_fd_sc_hd__xnor2_2 _27564_ (.A(_17705_),
    .B(_17715_),
    .Y(_17716_));
 sky130_fd_sc_hd__xnor2_2 _27565_ (.A(_17704_),
    .B(_17716_),
    .Y(_17717_));
 sky130_fd_sc_hd__and2_2 _27566_ (.A(_17483_),
    .B(_17487_),
    .X(_17718_));
 sky130_fd_sc_hd__xnor2_2 _27567_ (.A(_17717_),
    .B(_17718_),
    .Y(_17719_));
 sky130_fd_sc_hd__xnor2_2 _27568_ (.A(_17701_),
    .B(_17719_),
    .Y(_17720_));
 sky130_fd_sc_hd__and2_2 _27569_ (.A(_17491_),
    .B(_17493_),
    .X(_17721_));
 sky130_fd_sc_hd__xor2_2 _27570_ (.A(_17720_),
    .B(_17721_),
    .X(_17722_));
 sky130_fd_sc_hd__xnor2_2 _27571_ (.A(_17695_),
    .B(_17722_),
    .Y(_17723_));
 sky130_fd_sc_hd__nand2_2 _27572_ (.A(_17497_),
    .B(_17499_),
    .Y(_17724_));
 sky130_fd_sc_hd__xnor2_2 _27573_ (.A(_17723_),
    .B(_17724_),
    .Y(_17726_));
 sky130_fd_sc_hd__xor2_2 _27574_ (.A(_17682_),
    .B(_17726_),
    .X(_17727_));
 sky130_fd_sc_hd__nor2_2 _27575_ (.A(_17501_),
    .B(_17503_),
    .Y(_17728_));
 sky130_fd_sc_hd__xnor2_2 _27576_ (.A(_17727_),
    .B(_17728_),
    .Y(_17729_));
 sky130_fd_sc_hd__xnor2_2 _27577_ (.A(_17660_),
    .B(_17729_),
    .Y(_17730_));
 sky130_fd_sc_hd__a21bo_2 _27578_ (.A1(_17435_),
    .A2(_17509_),
    .B1_N(_17507_),
    .X(_17731_));
 sky130_fd_sc_hd__xor2_2 _27579_ (.A(_17730_),
    .B(_17731_),
    .X(_17732_));
 sky130_fd_sc_hd__xor2_2 _27580_ (.A(_17616_),
    .B(_17732_),
    .X(_17733_));
 sky130_fd_sc_hd__a21oi_2 _27581_ (.A1(_17381_),
    .A2(_17512_),
    .B1(_17511_),
    .Y(_17734_));
 sky130_fd_sc_hd__xor2_2 _27582_ (.A(_17733_),
    .B(_17734_),
    .X(_17735_));
 sky130_fd_sc_hd__xor2_2 _27583_ (.A(_17610_),
    .B(_17735_),
    .X(_17737_));
 sky130_fd_sc_hd__xor2_2 _27584_ (.A(_17609_),
    .B(_17737_),
    .X(_17738_));
 sky130_fd_sc_hd__xnor2_2 _27585_ (.A(_17608_),
    .B(_17738_),
    .Y(_17739_));
 sky130_fd_sc_hd__inv_2 _27586_ (.A(_17739_),
    .Y(_17740_));
 sky130_fd_sc_hd__nand2_2 _27587_ (.A(_17377_),
    .B(_17518_),
    .Y(_17741_));
 sky130_fd_sc_hd__o21ai_2 _27588_ (.A1(_17523_),
    .A2(_17519_),
    .B1(_17741_),
    .Y(_17742_));
 sky130_fd_sc_hd__a31o_2 _27589_ (.A1(_16900_),
    .A2(_17044_),
    .A3(_17520_),
    .B1(_17742_),
    .X(_17743_));
 sky130_fd_sc_hd__xnor2_2 _27590_ (.A(_17740_),
    .B(_17743_),
    .Y(_17744_));
 sky130_fd_sc_hd__inv_2 _27591_ (.A(_17157_),
    .Y(_17745_));
 sky130_fd_sc_hd__nor2_2 _27592_ (.A(_17745_),
    .B(_17370_),
    .Y(_17746_));
 sky130_fd_sc_hd__or2_2 _27593_ (.A(_17368_),
    .B(_17369_),
    .X(_17748_));
 sky130_fd_sc_hd__and3_2 _27594_ (.A(_17313_),
    .B(_17314_),
    .C(_17316_),
    .X(_17749_));
 sky130_fd_sc_hd__and2b_2 _27595_ (.A_N(_17277_),
    .B(_17276_),
    .X(_17750_));
 sky130_fd_sc_hd__and2_2 _27596_ (.A(_17270_),
    .B(_17278_),
    .X(_17751_));
 sky130_fd_sc_hd__or2b_2 _27597_ (.A(_17304_),
    .B_N(_17310_),
    .X(_17752_));
 sky130_fd_sc_hd__or2b_2 _27598_ (.A(_17303_),
    .B_N(_17311_),
    .X(_17753_));
 sky130_fd_sc_hd__and4_2 _27599_ (.A(iX[41]),
    .B(iX[42]),
    .C(iY[44]),
    .D(iY[45]),
    .X(_17754_));
 sky130_fd_sc_hd__a22oi_2 _27600_ (.A1(iX[42]),
    .A2(iY[44]),
    .B1(iY[45]),
    .B2(iX[41]),
    .Y(_17755_));
 sky130_fd_sc_hd__nor2_2 _27601_ (.A(_17754_),
    .B(_17755_),
    .Y(_17756_));
 sky130_fd_sc_hd__nand2_2 _27602_ (.A(iX[40]),
    .B(iY[46]),
    .Y(_17757_));
 sky130_fd_sc_hd__xnor2_2 _27603_ (.A(_17756_),
    .B(_17757_),
    .Y(_17759_));
 sky130_fd_sc_hd__and4_2 _27604_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[44]),
    .D(iX[45]),
    .X(_17760_));
 sky130_fd_sc_hd__a22oi_2 _27605_ (.A1(iY[42]),
    .A2(iX[44]),
    .B1(iX[45]),
    .B2(iY[41]),
    .Y(_17761_));
 sky130_fd_sc_hd__nor2_2 _27606_ (.A(_17760_),
    .B(_17761_),
    .Y(_17762_));
 sky130_fd_sc_hd__nand2_2 _27607_ (.A(iX[43]),
    .B(iY[43]),
    .Y(_17763_));
 sky130_fd_sc_hd__xnor2_2 _27608_ (.A(_17762_),
    .B(_17763_),
    .Y(_17764_));
 sky130_fd_sc_hd__o21ba_2 _27609_ (.A1(_17272_),
    .A2(_17274_),
    .B1_N(_17271_),
    .X(_17765_));
 sky130_fd_sc_hd__xnor2_2 _27610_ (.A(_17764_),
    .B(_17765_),
    .Y(_17766_));
 sky130_fd_sc_hd__and2_2 _27611_ (.A(_17759_),
    .B(_17766_),
    .X(_17767_));
 sky130_fd_sc_hd__nor2_2 _27612_ (.A(_17759_),
    .B(_17766_),
    .Y(_17768_));
 sky130_fd_sc_hd__or2_2 _27613_ (.A(_17767_),
    .B(_17768_),
    .X(_17770_));
 sky130_fd_sc_hd__a21o_2 _27614_ (.A1(_17752_),
    .A2(_17753_),
    .B1(_17770_),
    .X(_17771_));
 sky130_fd_sc_hd__nand3_2 _27615_ (.A(_17752_),
    .B(_17753_),
    .C(_17770_),
    .Y(_17772_));
 sky130_fd_sc_hd__o211ai_2 _27616_ (.A1(_17750_),
    .A2(_17751_),
    .B1(_17771_),
    .C1(_17772_),
    .Y(_17773_));
 sky130_fd_sc_hd__a211o_2 _27617_ (.A1(_17771_),
    .A2(_17772_),
    .B1(_17750_),
    .C1(_17751_),
    .X(_17774_));
 sky130_fd_sc_hd__or2b_2 _27618_ (.A(_17292_),
    .B_N(_17291_),
    .X(_17775_));
 sky130_fd_sc_hd__nand2_2 _27619_ (.A(_17293_),
    .B(_17299_),
    .Y(_17776_));
 sky130_fd_sc_hd__and4_2 _27620_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[51]),
    .D(iX[52]),
    .X(_17777_));
 sky130_fd_sc_hd__a22oi_2 _27621_ (.A1(iY[35]),
    .A2(iX[51]),
    .B1(iX[52]),
    .B2(iY[34]),
    .Y(_17778_));
 sky130_fd_sc_hd__nor2_2 _27622_ (.A(_17777_),
    .B(_17778_),
    .Y(_17779_));
 sky130_fd_sc_hd__nand2_2 _27623_ (.A(iY[33]),
    .B(iX[53]),
    .Y(_17781_));
 sky130_fd_sc_hd__xnor2_2 _27624_ (.A(_17779_),
    .B(_17781_),
    .Y(_17782_));
 sky130_fd_sc_hd__o21ba_2 _27625_ (.A1(_17288_),
    .A2(_17290_),
    .B1_N(_17287_),
    .X(_17783_));
 sky130_fd_sc_hd__xnor2_2 _27626_ (.A(_17782_),
    .B(_17783_),
    .Y(_17784_));
 sky130_fd_sc_hd__and4_2 _27627_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[50]),
    .D(iX[54]),
    .X(_17785_));
 sky130_fd_sc_hd__a22oi_2 _27628_ (.A1(iY[36]),
    .A2(iX[50]),
    .B1(iX[54]),
    .B2(iY[32]),
    .Y(_17786_));
 sky130_fd_sc_hd__nor2_2 _27629_ (.A(_17785_),
    .B(_17786_),
    .Y(_17787_));
 sky130_fd_sc_hd__nand2_2 _27630_ (.A(iY[37]),
    .B(iX[49]),
    .Y(_17788_));
 sky130_fd_sc_hd__xnor2_2 _27631_ (.A(_17787_),
    .B(_17788_),
    .Y(_17789_));
 sky130_fd_sc_hd__xnor2_2 _27632_ (.A(_17784_),
    .B(_17789_),
    .Y(_17790_));
 sky130_fd_sc_hd__a21o_2 _27633_ (.A1(_17775_),
    .A2(_17776_),
    .B1(_17790_),
    .X(_17792_));
 sky130_fd_sc_hd__nand3_2 _27634_ (.A(_17775_),
    .B(_17776_),
    .C(_17790_),
    .Y(_17793_));
 sky130_fd_sc_hd__o21ba_2 _27635_ (.A1(_17306_),
    .A2(_17309_),
    .B1_N(_17305_),
    .X(_17794_));
 sky130_fd_sc_hd__o21ba_2 _27636_ (.A1(_17295_),
    .A2(_17298_),
    .B1_N(_17294_),
    .X(_17795_));
 sky130_fd_sc_hd__and4_2 _27637_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[47]),
    .D(iX[48]),
    .X(_17796_));
 sky130_fd_sc_hd__a22oi_2 _27638_ (.A1(iY[39]),
    .A2(iX[47]),
    .B1(iX[48]),
    .B2(iY[38]),
    .Y(_17797_));
 sky130_fd_sc_hd__nor2_2 _27639_ (.A(_17796_),
    .B(_17797_),
    .Y(_17798_));
 sky130_fd_sc_hd__nand2_2 _27640_ (.A(iY[40]),
    .B(iX[46]),
    .Y(_17799_));
 sky130_fd_sc_hd__xnor2_2 _27641_ (.A(_17798_),
    .B(_17799_),
    .Y(_17800_));
 sky130_fd_sc_hd__xnor2_2 _27642_ (.A(_17795_),
    .B(_17800_),
    .Y(_17801_));
 sky130_fd_sc_hd__xnor2_2 _27643_ (.A(_17794_),
    .B(_17801_),
    .Y(_17803_));
 sky130_fd_sc_hd__nand3_2 _27644_ (.A(_17792_),
    .B(_17793_),
    .C(_17803_),
    .Y(_17804_));
 sky130_fd_sc_hd__a21o_2 _27645_ (.A1(_17792_),
    .A2(_17793_),
    .B1(_17803_),
    .X(_17805_));
 sky130_fd_sc_hd__nand2_2 _27646_ (.A(_17804_),
    .B(_17805_),
    .Y(_17806_));
 sky130_fd_sc_hd__nand2_2 _27647_ (.A(_17301_),
    .B(_17313_),
    .Y(_17807_));
 sky130_fd_sc_hd__xnor2_2 _27648_ (.A(_17806_),
    .B(_17807_),
    .Y(_17808_));
 sky130_fd_sc_hd__a21o_2 _27649_ (.A1(_17773_),
    .A2(_17774_),
    .B1(_17808_),
    .X(_17809_));
 sky130_fd_sc_hd__nand3_2 _27650_ (.A(_17808_),
    .B(_17773_),
    .C(_17774_),
    .Y(_17810_));
 sky130_fd_sc_hd__o211a_2 _27651_ (.A1(_17749_),
    .A2(_17320_),
    .B1(_17809_),
    .C1(_17810_),
    .X(_17811_));
 sky130_fd_sc_hd__a211oi_2 _27652_ (.A1(_17809_),
    .A2(_17810_),
    .B1(_17749_),
    .C1(_17320_),
    .Y(_17812_));
 sky130_fd_sc_hd__inv_2 _27653_ (.A(_17347_),
    .Y(_17814_));
 sky130_fd_sc_hd__a22oi_2 _27654_ (.A1(iX[33]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[32]),
    .Y(_17815_));
 sky130_fd_sc_hd__and4_2 _27655_ (.A(iX[33]),
    .B(iX[32]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_17816_));
 sky130_fd_sc_hd__or2_2 _27656_ (.A(_17815_),
    .B(_17816_),
    .X(_17817_));
 sky130_fd_sc_hd__and4_2 _27657_ (.A(iX[35]),
    .B(iX[36]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_17818_));
 sky130_fd_sc_hd__a22o_2 _27658_ (.A1(iX[36]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[35]),
    .X(_17819_));
 sky130_fd_sc_hd__and2b_2 _27659_ (.A_N(_17818_),
    .B(_17819_),
    .X(_17820_));
 sky130_fd_sc_hd__nand2_2 _27660_ (.A(iX[34]),
    .B(iY[52]),
    .Y(_17821_));
 sky130_fd_sc_hd__xnor2_2 _27661_ (.A(_17820_),
    .B(_17821_),
    .Y(_17822_));
 sky130_fd_sc_hd__o21ba_2 _27662_ (.A1(_17326_),
    .A2(_17328_),
    .B1_N(_17325_),
    .X(_17823_));
 sky130_fd_sc_hd__xnor2_2 _27663_ (.A(_17822_),
    .B(_17823_),
    .Y(_17825_));
 sky130_fd_sc_hd__xnor2_2 _27664_ (.A(_17817_),
    .B(_17825_),
    .Y(_17826_));
 sky130_fd_sc_hd__or2b_2 _27665_ (.A(_17336_),
    .B_N(_17342_),
    .X(_17827_));
 sky130_fd_sc_hd__a31o_2 _27666_ (.A1(iX[36]),
    .A2(iY[49]),
    .A3(_17339_),
    .B1(_17337_),
    .X(_17828_));
 sky130_fd_sc_hd__o21ba_2 _27667_ (.A1(_17267_),
    .A2(_17269_),
    .B1_N(_17266_),
    .X(_17829_));
 sky130_fd_sc_hd__and4_2 _27668_ (.A(iX[38]),
    .B(iX[39]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_17830_));
 sky130_fd_sc_hd__a22oi_2 _27669_ (.A1(iX[39]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[38]),
    .Y(_17831_));
 sky130_fd_sc_hd__nor2_2 _27670_ (.A(_17830_),
    .B(_17831_),
    .Y(_17832_));
 sky130_fd_sc_hd__nand2_2 _27671_ (.A(iX[37]),
    .B(iY[49]),
    .Y(_17833_));
 sky130_fd_sc_hd__xnor2_2 _27672_ (.A(_17832_),
    .B(_17833_),
    .Y(_17834_));
 sky130_fd_sc_hd__xnor2_2 _27673_ (.A(_17829_),
    .B(_17834_),
    .Y(_17835_));
 sky130_fd_sc_hd__xnor2_2 _27674_ (.A(_17828_),
    .B(_17835_),
    .Y(_17836_));
 sky130_fd_sc_hd__a21o_2 _27675_ (.A1(_17827_),
    .A2(_17344_),
    .B1(_17836_),
    .X(_17837_));
 sky130_fd_sc_hd__nand3_2 _27676_ (.A(_17827_),
    .B(_17344_),
    .C(_17836_),
    .Y(_17838_));
 sky130_fd_sc_hd__and3_2 _27677_ (.A(_17826_),
    .B(_17837_),
    .C(_17838_),
    .X(_17839_));
 sky130_fd_sc_hd__a21oi_2 _27678_ (.A1(_17837_),
    .A2(_17838_),
    .B1(_17826_),
    .Y(_17840_));
 sky130_fd_sc_hd__a211o_2 _27679_ (.A1(_17280_),
    .A2(_17282_),
    .B1(_17839_),
    .C1(_17840_),
    .X(_17841_));
 sky130_fd_sc_hd__inv_2 _27680_ (.A(_17841_),
    .Y(_17842_));
 sky130_fd_sc_hd__o211a_2 _27681_ (.A1(_17839_),
    .A2(_17840_),
    .B1(_17280_),
    .C1(_17282_),
    .X(_17843_));
 sky130_fd_sc_hd__a211o_2 _27682_ (.A1(_17814_),
    .A2(_17349_),
    .B1(_17842_),
    .C1(_17843_),
    .X(_17844_));
 sky130_fd_sc_hd__inv_2 _27683_ (.A(_17844_),
    .Y(_17846_));
 sky130_fd_sc_hd__o211a_2 _27684_ (.A1(_17842_),
    .A2(_17843_),
    .B1(_17814_),
    .C1(_17349_),
    .X(_17847_));
 sky130_fd_sc_hd__nor4_2 _27685_ (.A(_17811_),
    .B(_17812_),
    .C(_17846_),
    .D(_17847_),
    .Y(_17848_));
 sky130_fd_sc_hd__o22a_2 _27686_ (.A1(_17811_),
    .A2(_17812_),
    .B1(_17846_),
    .B2(_17847_),
    .X(_17849_));
 sky130_fd_sc_hd__a211o_2 _27687_ (.A1(_17322_),
    .A2(_17358_),
    .B1(_17848_),
    .C1(_17849_),
    .X(_17850_));
 sky130_fd_sc_hd__o211ai_2 _27688_ (.A1(_17848_),
    .A2(_17849_),
    .B1(_17322_),
    .C1(_17358_),
    .Y(_17851_));
 sky130_fd_sc_hd__and2b_2 _27689_ (.A_N(_17331_),
    .B(_17329_),
    .X(_17852_));
 sky130_fd_sc_hd__a31oi_2 _27690_ (.A1(iX[32]),
    .A2(iY[53]),
    .A3(_17332_),
    .B1(_17852_),
    .Y(_17853_));
 sky130_fd_sc_hd__o21ba_2 _27691_ (.A1(_17353_),
    .A2(_17355_),
    .B1_N(_17853_),
    .X(_17854_));
 sky130_fd_sc_hd__or3b_2 _27692_ (.A(_17353_),
    .B(_17355_),
    .C_N(_17853_),
    .X(_17855_));
 sky130_fd_sc_hd__and2b_2 _27693_ (.A_N(_17854_),
    .B(_17855_),
    .X(_17857_));
 sky130_fd_sc_hd__and3_2 _27694_ (.A(_17850_),
    .B(_17851_),
    .C(_17857_),
    .X(_17858_));
 sky130_fd_sc_hd__a21oi_2 _27695_ (.A1(_17850_),
    .A2(_17851_),
    .B1(_17857_),
    .Y(_17859_));
 sky130_fd_sc_hd__nor2_2 _27696_ (.A(_17858_),
    .B(_17859_),
    .Y(_17860_));
 sky130_fd_sc_hd__a21bo_2 _27697_ (.A1(_17361_),
    .A2(_17365_),
    .B1_N(_17360_),
    .X(_17861_));
 sky130_fd_sc_hd__xnor2_2 _27698_ (.A(_17860_),
    .B(_17861_),
    .Y(_17862_));
 sky130_fd_sc_hd__xnor2_2 _27699_ (.A(_17362_),
    .B(_17862_),
    .Y(_17863_));
 sky130_fd_sc_hd__xor2_2 _27700_ (.A(_17748_),
    .B(_17863_),
    .X(_17864_));
 sky130_fd_sc_hd__xnor2_2 _27701_ (.A(_17746_),
    .B(_17864_),
    .Y(_17865_));
 sky130_fd_sc_hd__and2b_2 _27702_ (.A_N(_17159_),
    .B(_17371_),
    .X(_17866_));
 sky130_fd_sc_hd__nor2_2 _27703_ (.A(_17866_),
    .B(_17375_),
    .Y(_17868_));
 sky130_fd_sc_hd__xor2_2 _27704_ (.A(_17865_),
    .B(_17868_),
    .X(_17869_));
 sky130_fd_sc_hd__xor2_2 _27705_ (.A(_17744_),
    .B(_17869_),
    .X(_17870_));
 sky130_fd_sc_hd__xor2_2 _27706_ (.A(oO[22]),
    .B(_17870_),
    .X(_17871_));
 sky130_fd_sc_hd__a21oi_2 _27707_ (.A1(_17606_),
    .A2(_17607_),
    .B1(_17871_),
    .Y(_17872_));
 sky130_fd_sc_hd__inv_2 _27708_ (.A(_17872_),
    .Y(_17873_));
 sky130_fd_sc_hd__nand3_2 _27709_ (.A(_17606_),
    .B(_17607_),
    .C(_17871_),
    .Y(_17874_));
 sky130_fd_sc_hd__nand2_2 _27710_ (.A(_17873_),
    .B(_17874_),
    .Y(_17875_));
 sky130_fd_sc_hd__or2b_2 _27711_ (.A(_17180_),
    .B_N(_17530_),
    .X(_17876_));
 sky130_fd_sc_hd__a31o_2 _27712_ (.A1(_16891_),
    .A2(_16730_),
    .A3(_16731_),
    .B1(_17876_),
    .X(_17877_));
 sky130_fd_sc_hd__and2b_2 _27713_ (.A_N(_17529_),
    .B(_17527_),
    .X(_17879_));
 sky130_fd_sc_hd__a21oi_2 _27714_ (.A1(_17531_),
    .A2(_17530_),
    .B1(_17879_),
    .Y(_17880_));
 sky130_fd_sc_hd__and2_2 _27715_ (.A(_17877_),
    .B(_17880_),
    .X(_17881_));
 sky130_fd_sc_hd__xnor2_2 _27716_ (.A(_17875_),
    .B(_17881_),
    .Y(_17882_));
 sky130_fd_sc_hd__nor2_2 _27717_ (.A(_17605_),
    .B(_17882_),
    .Y(_17883_));
 sky130_fd_sc_hd__and2_2 _27718_ (.A(_17605_),
    .B(_17882_),
    .X(_17884_));
 sky130_fd_sc_hd__nor2_2 _27719_ (.A(_17883_),
    .B(_17884_),
    .Y(_17885_));
 sky130_fd_sc_hd__nand2_2 _27720_ (.A(_17259_),
    .B(_17533_),
    .Y(_17886_));
 sky130_fd_sc_hd__o21ai_2 _27721_ (.A1(_17537_),
    .A2(_17535_),
    .B1(_17886_),
    .Y(_17887_));
 sky130_fd_sc_hd__a21boi_2 _27722_ (.A1(_17538_),
    .A2(_17536_),
    .B1_N(_17887_),
    .Y(_17888_));
 sky130_fd_sc_hd__xnor2_2 _27723_ (.A(_17885_),
    .B(_17888_),
    .Y(oO[54]));
 sky130_fd_sc_hd__o21ai_2 _27724_ (.A1(_17541_),
    .A2(_17587_),
    .B1(_17585_),
    .Y(_17890_));
 sky130_fd_sc_hd__and3_2 _27725_ (.A(iY[24]),
    .B(iX[31]),
    .C(_17543_),
    .X(_17891_));
 sky130_fd_sc_hd__a21o_2 _27726_ (.A1(iY[24]),
    .A2(iX[31]),
    .B1(_17543_),
    .X(_17892_));
 sky130_fd_sc_hd__and4b_2 _27727_ (.A_N(_17891_),
    .B(iX[29]),
    .C(iY[26]),
    .D(_17892_),
    .X(_17893_));
 sky130_fd_sc_hd__inv_2 _27728_ (.A(_17892_),
    .Y(_17894_));
 sky130_fd_sc_hd__o2bb2a_2 _27729_ (.A1_N(iY[26]),
    .A2_N(iX[29]),
    .B1(_17894_),
    .B2(_17891_),
    .X(_17895_));
 sky130_fd_sc_hd__nor2_2 _27730_ (.A(_17893_),
    .B(_17895_),
    .Y(_17896_));
 sky130_fd_sc_hd__or2_2 _27731_ (.A(_17544_),
    .B(_17546_),
    .X(_17897_));
 sky130_fd_sc_hd__xnor2_2 _27732_ (.A(_17896_),
    .B(_17897_),
    .Y(_17898_));
 sky130_fd_sc_hd__a21oi_2 _27733_ (.A1(_17195_),
    .A2(_17548_),
    .B1(_17552_),
    .Y(_17900_));
 sky130_fd_sc_hd__nor2_2 _27734_ (.A(_17898_),
    .B(_17900_),
    .Y(_17901_));
 sky130_fd_sc_hd__and2_2 _27735_ (.A(_17898_),
    .B(_17900_),
    .X(_17902_));
 sky130_fd_sc_hd__nor2_2 _27736_ (.A(_17901_),
    .B(_17902_),
    .Y(_17903_));
 sky130_fd_sc_hd__or2_2 _27737_ (.A(_17555_),
    .B(_17903_),
    .X(_17904_));
 sky130_fd_sc_hd__nand2_2 _27738_ (.A(_17555_),
    .B(_17903_),
    .Y(_17905_));
 sky130_fd_sc_hd__and2_2 _27739_ (.A(_17904_),
    .B(_17905_),
    .X(_17906_));
 sky130_fd_sc_hd__or2b_2 _27740_ (.A(_17566_),
    .B_N(_17565_),
    .X(_17907_));
 sky130_fd_sc_hd__and4_2 _27741_ (.A(iX[27]),
    .B(iY[27]),
    .C(iX[28]),
    .D(iY[28]),
    .X(_17908_));
 sky130_fd_sc_hd__a22oi_2 _27742_ (.A1(iY[27]),
    .A2(iX[28]),
    .B1(iY[28]),
    .B2(iX[27]),
    .Y(_17909_));
 sky130_fd_sc_hd__nor2_2 _27743_ (.A(_17908_),
    .B(_17909_),
    .Y(_17911_));
 sky130_fd_sc_hd__nand2_2 _27744_ (.A(iX[26]),
    .B(iY[29]),
    .Y(_17912_));
 sky130_fd_sc_hd__xnor2_2 _27745_ (.A(_17911_),
    .B(_17912_),
    .Y(_17913_));
 sky130_fd_sc_hd__o21ba_2 _27746_ (.A1(_17562_),
    .A2(_17564_),
    .B1_N(_17561_),
    .X(_17914_));
 sky130_fd_sc_hd__xnor2_2 _27747_ (.A(_17913_),
    .B(_17914_),
    .Y(_17915_));
 sky130_fd_sc_hd__nand3_2 _27748_ (.A(iX[25]),
    .B(iY[30]),
    .C(_17915_),
    .Y(_17916_));
 sky130_fd_sc_hd__a21o_2 _27749_ (.A1(iX[25]),
    .A2(iY[30]),
    .B1(_17915_),
    .X(_17917_));
 sky130_fd_sc_hd__nand2_2 _27750_ (.A(_17916_),
    .B(_17917_),
    .Y(_17918_));
 sky130_fd_sc_hd__a21oi_2 _27751_ (.A1(_17907_),
    .A2(_17568_),
    .B1(_17918_),
    .Y(_17919_));
 sky130_fd_sc_hd__and3_2 _27752_ (.A(_17907_),
    .B(_17568_),
    .C(_17918_),
    .X(_17920_));
 sky130_fd_sc_hd__nor2_2 _27753_ (.A(_17919_),
    .B(_17920_),
    .Y(_17922_));
 sky130_fd_sc_hd__nand2_2 _27754_ (.A(iX[24]),
    .B(iY[31]),
    .Y(_17923_));
 sky130_fd_sc_hd__xnor2_2 _27755_ (.A(_17922_),
    .B(_17923_),
    .Y(_17924_));
 sky130_fd_sc_hd__or2_2 _27756_ (.A(_17906_),
    .B(_17924_),
    .X(_17925_));
 sky130_fd_sc_hd__nand2_2 _27757_ (.A(_17906_),
    .B(_17924_),
    .Y(_17926_));
 sky130_fd_sc_hd__a21bo_2 _27758_ (.A1(_17558_),
    .A2(_17576_),
    .B1_N(_17557_),
    .X(_17927_));
 sky130_fd_sc_hd__and3_2 _27759_ (.A(_17925_),
    .B(_17926_),
    .C(_17927_),
    .X(_17928_));
 sky130_fd_sc_hd__a21oi_2 _27760_ (.A1(_17925_),
    .A2(_17926_),
    .B1(_17927_),
    .Y(_17929_));
 sky130_fd_sc_hd__nor2_2 _27761_ (.A(_17928_),
    .B(_17929_),
    .Y(_17930_));
 sky130_fd_sc_hd__o21ai_2 _27762_ (.A1(_17542_),
    .A2(_17583_),
    .B1(_17580_),
    .Y(_17931_));
 sky130_fd_sc_hd__xor2_2 _27763_ (.A(_17930_),
    .B(_17931_),
    .X(_17933_));
 sky130_fd_sc_hd__xnor2_2 _27764_ (.A(_17890_),
    .B(_17933_),
    .Y(_17934_));
 sky130_fd_sc_hd__o21ba_2 _27765_ (.A1(_17573_),
    .A2(_17575_),
    .B1_N(_17572_),
    .X(_17935_));
 sky130_fd_sc_hd__nor2_2 _27766_ (.A(_17934_),
    .B(_17935_),
    .Y(_17936_));
 sky130_fd_sc_hd__and2_2 _27767_ (.A(_17934_),
    .B(_17935_),
    .X(_17937_));
 sky130_fd_sc_hd__or2_2 _27768_ (.A(_17936_),
    .B(_17937_),
    .X(_17938_));
 sky130_fd_sc_hd__and3_2 _27769_ (.A(_17591_),
    .B(_17596_),
    .C(_17938_),
    .X(_17939_));
 sky130_fd_sc_hd__a21o_2 _27770_ (.A1(_17591_),
    .A2(_17596_),
    .B1(_17938_),
    .X(_17940_));
 sky130_fd_sc_hd__or2b_2 _27771_ (.A(_17939_),
    .B_N(_17940_),
    .X(_17941_));
 sky130_fd_sc_hd__o21a_2 _27772_ (.A1(_17602_),
    .A2(_17603_),
    .B1(_17600_),
    .X(_17942_));
 sky130_fd_sc_hd__xnor2_2 _27773_ (.A(_17941_),
    .B(_17942_),
    .Y(_17944_));
 sky130_fd_sc_hd__o21ai_2 _27774_ (.A1(_17875_),
    .A2(_17881_),
    .B1(_17873_),
    .Y(_17945_));
 sky130_fd_sc_hd__or2_2 _27775_ (.A(_17744_),
    .B(_17869_),
    .X(_17946_));
 sky130_fd_sc_hd__or2b_2 _27776_ (.A(oO[22]),
    .B_N(_17870_),
    .X(_17947_));
 sky130_fd_sc_hd__or2_2 _27777_ (.A(_17748_),
    .B(_17863_),
    .X(_17948_));
 sky130_fd_sc_hd__or2b_2 _27778_ (.A(_17806_),
    .B_N(_17807_),
    .X(_17949_));
 sky130_fd_sc_hd__or2b_2 _27779_ (.A(_17783_),
    .B_N(_17782_),
    .X(_17950_));
 sky130_fd_sc_hd__nand2_2 _27780_ (.A(_17784_),
    .B(_17789_),
    .Y(_17951_));
 sky130_fd_sc_hd__and4_2 _27781_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[52]),
    .D(iX[53]),
    .X(_17952_));
 sky130_fd_sc_hd__a22oi_2 _27782_ (.A1(iY[35]),
    .A2(iX[52]),
    .B1(iX[53]),
    .B2(iY[34]),
    .Y(_17953_));
 sky130_fd_sc_hd__nor2_2 _27783_ (.A(_17952_),
    .B(_17953_),
    .Y(_17955_));
 sky130_fd_sc_hd__nand2_2 _27784_ (.A(iY[33]),
    .B(iX[54]),
    .Y(_17956_));
 sky130_fd_sc_hd__xnor2_2 _27785_ (.A(_17955_),
    .B(_17956_),
    .Y(_17957_));
 sky130_fd_sc_hd__o21ba_2 _27786_ (.A1(_17778_),
    .A2(_17781_),
    .B1_N(_17777_),
    .X(_17958_));
 sky130_fd_sc_hd__xnor2_2 _27787_ (.A(_17957_),
    .B(_17958_),
    .Y(_17959_));
 sky130_fd_sc_hd__and4_2 _27788_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[51]),
    .D(iX[55]),
    .X(_17960_));
 sky130_fd_sc_hd__a22oi_2 _27789_ (.A1(iY[36]),
    .A2(iX[51]),
    .B1(iX[55]),
    .B2(iY[32]),
    .Y(_17961_));
 sky130_fd_sc_hd__nor2_2 _27790_ (.A(_17960_),
    .B(_17961_),
    .Y(_17962_));
 sky130_fd_sc_hd__nand2_2 _27791_ (.A(iY[37]),
    .B(iX[50]),
    .Y(_17963_));
 sky130_fd_sc_hd__xnor2_2 _27792_ (.A(_17962_),
    .B(_17963_),
    .Y(_17964_));
 sky130_fd_sc_hd__xnor2_2 _27793_ (.A(_17959_),
    .B(_17964_),
    .Y(_17966_));
 sky130_fd_sc_hd__a21o_2 _27794_ (.A1(_17950_),
    .A2(_17951_),
    .B1(_17966_),
    .X(_17967_));
 sky130_fd_sc_hd__nand3_2 _27795_ (.A(_17950_),
    .B(_17951_),
    .C(_17966_),
    .Y(_17968_));
 sky130_fd_sc_hd__o21ba_2 _27796_ (.A1(_17797_),
    .A2(_17799_),
    .B1_N(_17796_),
    .X(_17969_));
 sky130_fd_sc_hd__o21ba_2 _27797_ (.A1(_17786_),
    .A2(_17788_),
    .B1_N(_17785_),
    .X(_17970_));
 sky130_fd_sc_hd__and4_2 _27798_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[48]),
    .D(iX[49]),
    .X(_17971_));
 sky130_fd_sc_hd__a22oi_2 _27799_ (.A1(iY[39]),
    .A2(iX[48]),
    .B1(iX[49]),
    .B2(iY[38]),
    .Y(_17972_));
 sky130_fd_sc_hd__nor2_2 _27800_ (.A(_17971_),
    .B(_17972_),
    .Y(_17973_));
 sky130_fd_sc_hd__nand2_2 _27801_ (.A(iY[40]),
    .B(iX[47]),
    .Y(_17974_));
 sky130_fd_sc_hd__xnor2_2 _27802_ (.A(_17973_),
    .B(_17974_),
    .Y(_17975_));
 sky130_fd_sc_hd__xnor2_2 _27803_ (.A(_17970_),
    .B(_17975_),
    .Y(_17977_));
 sky130_fd_sc_hd__xnor2_2 _27804_ (.A(_17969_),
    .B(_17977_),
    .Y(_17978_));
 sky130_fd_sc_hd__nand3_2 _27805_ (.A(_17967_),
    .B(_17968_),
    .C(_17978_),
    .Y(_17979_));
 sky130_fd_sc_hd__a21o_2 _27806_ (.A1(_17967_),
    .A2(_17968_),
    .B1(_17978_),
    .X(_17980_));
 sky130_fd_sc_hd__nand2_2 _27807_ (.A(_17979_),
    .B(_17980_),
    .Y(_17981_));
 sky130_fd_sc_hd__nand2_2 _27808_ (.A(_17792_),
    .B(_17804_),
    .Y(_17982_));
 sky130_fd_sc_hd__xnor2_2 _27809_ (.A(_17981_),
    .B(_17982_),
    .Y(_17983_));
 sky130_fd_sc_hd__and2b_2 _27810_ (.A_N(_17765_),
    .B(_17764_),
    .X(_17984_));
 sky130_fd_sc_hd__or2b_2 _27811_ (.A(_17795_),
    .B_N(_17800_),
    .X(_17985_));
 sky130_fd_sc_hd__or2b_2 _27812_ (.A(_17794_),
    .B_N(_17801_),
    .X(_17986_));
 sky130_fd_sc_hd__and4_2 _27813_ (.A(iX[42]),
    .B(iX[43]),
    .C(iY[44]),
    .D(iY[45]),
    .X(_17988_));
 sky130_fd_sc_hd__a22oi_2 _27814_ (.A1(iX[43]),
    .A2(iY[44]),
    .B1(iY[45]),
    .B2(iX[42]),
    .Y(_17989_));
 sky130_fd_sc_hd__nor2_2 _27815_ (.A(_17988_),
    .B(_17989_),
    .Y(_17990_));
 sky130_fd_sc_hd__nand2_2 _27816_ (.A(iX[41]),
    .B(iY[46]),
    .Y(_17991_));
 sky130_fd_sc_hd__xnor2_2 _27817_ (.A(_17990_),
    .B(_17991_),
    .Y(_17992_));
 sky130_fd_sc_hd__and4_2 _27818_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[45]),
    .D(iX[46]),
    .X(_17993_));
 sky130_fd_sc_hd__a22oi_2 _27819_ (.A1(iY[42]),
    .A2(iX[45]),
    .B1(iX[46]),
    .B2(iY[41]),
    .Y(_17994_));
 sky130_fd_sc_hd__and4bb_2 _27820_ (.A_N(_17993_),
    .B_N(_17994_),
    .C(iY[43]),
    .D(iX[44]),
    .X(_17995_));
 sky130_fd_sc_hd__o2bb2a_2 _27821_ (.A1_N(iY[43]),
    .A2_N(iX[44]),
    .B1(_17993_),
    .B2(_17994_),
    .X(_17996_));
 sky130_fd_sc_hd__nor2_2 _27822_ (.A(_17995_),
    .B(_17996_),
    .Y(_17997_));
 sky130_fd_sc_hd__o21ba_2 _27823_ (.A1(_17761_),
    .A2(_17763_),
    .B1_N(_17760_),
    .X(_17999_));
 sky130_fd_sc_hd__xnor2_2 _27824_ (.A(_17997_),
    .B(_17999_),
    .Y(_18000_));
 sky130_fd_sc_hd__and2_2 _27825_ (.A(_17992_),
    .B(_18000_),
    .X(_18001_));
 sky130_fd_sc_hd__nor2_2 _27826_ (.A(_17992_),
    .B(_18000_),
    .Y(_18002_));
 sky130_fd_sc_hd__or2_2 _27827_ (.A(_18001_),
    .B(_18002_),
    .X(_18003_));
 sky130_fd_sc_hd__a21o_2 _27828_ (.A1(_17985_),
    .A2(_17986_),
    .B1(_18003_),
    .X(_18004_));
 sky130_fd_sc_hd__nand3_2 _27829_ (.A(_17985_),
    .B(_17986_),
    .C(_18003_),
    .Y(_18005_));
 sky130_fd_sc_hd__o211ai_2 _27830_ (.A1(_17984_),
    .A2(_17767_),
    .B1(_18004_),
    .C1(_18005_),
    .Y(_18006_));
 sky130_fd_sc_hd__a211o_2 _27831_ (.A1(_18004_),
    .A2(_18005_),
    .B1(_17984_),
    .C1(_17767_),
    .X(_18007_));
 sky130_fd_sc_hd__and3_2 _27832_ (.A(_17983_),
    .B(_18006_),
    .C(_18007_),
    .X(_18008_));
 sky130_fd_sc_hd__a21oi_2 _27833_ (.A1(_18006_),
    .A2(_18007_),
    .B1(_17983_),
    .Y(_18010_));
 sky130_fd_sc_hd__a211o_2 _27834_ (.A1(_17949_),
    .A2(_17810_),
    .B1(_18008_),
    .C1(_18010_),
    .X(_18011_));
 sky130_fd_sc_hd__o211ai_2 _27835_ (.A1(_18008_),
    .A2(_18010_),
    .B1(_17949_),
    .C1(_17810_),
    .Y(_18012_));
 sky130_fd_sc_hd__inv_2 _27836_ (.A(_17839_),
    .Y(_18013_));
 sky130_fd_sc_hd__and4_2 _27837_ (.A(iX[33]),
    .B(iX[34]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_18014_));
 sky130_fd_sc_hd__a22o_2 _27838_ (.A1(iX[34]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[33]),
    .X(_18015_));
 sky130_fd_sc_hd__and2b_2 _27839_ (.A_N(_18014_),
    .B(_18015_),
    .X(_18016_));
 sky130_fd_sc_hd__nand2_2 _27840_ (.A(iX[32]),
    .B(iY[55]),
    .Y(_18017_));
 sky130_fd_sc_hd__xnor2_2 _27841_ (.A(_18016_),
    .B(_18017_),
    .Y(_18018_));
 sky130_fd_sc_hd__and4_2 _27842_ (.A(iX[36]),
    .B(iX[37]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_18019_));
 sky130_fd_sc_hd__a22o_2 _27843_ (.A1(iX[37]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[36]),
    .X(_18021_));
 sky130_fd_sc_hd__and2b_2 _27844_ (.A_N(_18019_),
    .B(_18021_),
    .X(_18022_));
 sky130_fd_sc_hd__nand2_2 _27845_ (.A(iX[35]),
    .B(iY[52]),
    .Y(_18023_));
 sky130_fd_sc_hd__xnor2_2 _27846_ (.A(_18022_),
    .B(_18023_),
    .Y(_18024_));
 sky130_fd_sc_hd__a31o_2 _27847_ (.A1(iX[34]),
    .A2(iY[52]),
    .A3(_17819_),
    .B1(_17818_),
    .X(_18025_));
 sky130_fd_sc_hd__xor2_2 _27848_ (.A(_18024_),
    .B(_18025_),
    .X(_18026_));
 sky130_fd_sc_hd__and2_2 _27849_ (.A(_18018_),
    .B(_18026_),
    .X(_18027_));
 sky130_fd_sc_hd__nor2_2 _27850_ (.A(_18018_),
    .B(_18026_),
    .Y(_18028_));
 sky130_fd_sc_hd__or2_2 _27851_ (.A(_18027_),
    .B(_18028_),
    .X(_18029_));
 sky130_fd_sc_hd__or2b_2 _27852_ (.A(_17829_),
    .B_N(_17834_),
    .X(_18030_));
 sky130_fd_sc_hd__nand2_2 _27853_ (.A(_17828_),
    .B(_17835_),
    .Y(_18032_));
 sky130_fd_sc_hd__a31o_2 _27854_ (.A1(iX[37]),
    .A2(iY[49]),
    .A3(_17832_),
    .B1(_17830_),
    .X(_18033_));
 sky130_fd_sc_hd__o21ba_2 _27855_ (.A1(_17755_),
    .A2(_17757_),
    .B1_N(_17754_),
    .X(_18034_));
 sky130_fd_sc_hd__and4_2 _27856_ (.A(iX[39]),
    .B(iX[40]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_18035_));
 sky130_fd_sc_hd__a22oi_2 _27857_ (.A1(iX[40]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[39]),
    .Y(_18036_));
 sky130_fd_sc_hd__and4bb_2 _27858_ (.A_N(_18035_),
    .B_N(_18036_),
    .C(iX[38]),
    .D(iY[49]),
    .X(_18037_));
 sky130_fd_sc_hd__o2bb2a_2 _27859_ (.A1_N(iX[38]),
    .A2_N(iY[49]),
    .B1(_18035_),
    .B2(_18036_),
    .X(_18038_));
 sky130_fd_sc_hd__nor2_2 _27860_ (.A(_18037_),
    .B(_18038_),
    .Y(_18039_));
 sky130_fd_sc_hd__xnor2_2 _27861_ (.A(_18034_),
    .B(_18039_),
    .Y(_18040_));
 sky130_fd_sc_hd__xnor2_2 _27862_ (.A(_18033_),
    .B(_18040_),
    .Y(_18041_));
 sky130_fd_sc_hd__a21oi_2 _27863_ (.A1(_18030_),
    .A2(_18032_),
    .B1(_18041_),
    .Y(_18043_));
 sky130_fd_sc_hd__and3_2 _27864_ (.A(_18030_),
    .B(_18032_),
    .C(_18041_),
    .X(_18044_));
 sky130_fd_sc_hd__or3_2 _27865_ (.A(_18029_),
    .B(_18043_),
    .C(_18044_),
    .X(_18045_));
 sky130_fd_sc_hd__o21ai_2 _27866_ (.A1(_18043_),
    .A2(_18044_),
    .B1(_18029_),
    .Y(_18046_));
 sky130_fd_sc_hd__nand2_2 _27867_ (.A(_18045_),
    .B(_18046_),
    .Y(_18047_));
 sky130_fd_sc_hd__a21oi_2 _27868_ (.A1(_17771_),
    .A2(_17773_),
    .B1(_18047_),
    .Y(_18048_));
 sky130_fd_sc_hd__and3_2 _27869_ (.A(_17771_),
    .B(_17773_),
    .C(_18047_),
    .X(_18049_));
 sky130_fd_sc_hd__a211oi_2 _27870_ (.A1(_17837_),
    .A2(_18013_),
    .B1(_18048_),
    .C1(_18049_),
    .Y(_18050_));
 sky130_fd_sc_hd__o211a_2 _27871_ (.A1(_18048_),
    .A2(_18049_),
    .B1(_17837_),
    .C1(_18013_),
    .X(_18051_));
 sky130_fd_sc_hd__nor2_2 _27872_ (.A(_18050_),
    .B(_18051_),
    .Y(_18052_));
 sky130_fd_sc_hd__and3_2 _27873_ (.A(_18011_),
    .B(_18012_),
    .C(_18052_),
    .X(_18054_));
 sky130_fd_sc_hd__a21oi_2 _27874_ (.A1(_18011_),
    .A2(_18012_),
    .B1(_18052_),
    .Y(_18055_));
 sky130_fd_sc_hd__nor2_2 _27875_ (.A(_18054_),
    .B(_18055_),
    .Y(_18056_));
 sky130_fd_sc_hd__nor2_2 _27876_ (.A(_17811_),
    .B(_17848_),
    .Y(_18057_));
 sky130_fd_sc_hd__xnor2_2 _27877_ (.A(_18056_),
    .B(_18057_),
    .Y(_18058_));
 sky130_fd_sc_hd__nand2_2 _27878_ (.A(_17841_),
    .B(_17844_),
    .Y(_18059_));
 sky130_fd_sc_hd__inv_2 _27879_ (.A(_17825_),
    .Y(_18060_));
 sky130_fd_sc_hd__and2b_2 _27880_ (.A_N(_17823_),
    .B(_17822_),
    .X(_18061_));
 sky130_fd_sc_hd__nand2_2 _27881_ (.A(_17816_),
    .B(_18061_),
    .Y(_18062_));
 sky130_fd_sc_hd__or2_2 _27882_ (.A(_17816_),
    .B(_18061_),
    .X(_18063_));
 sky130_fd_sc_hd__a2bb2o_2 _27883_ (.A1_N(_17817_),
    .A2_N(_18060_),
    .B1(_18062_),
    .B2(_18063_),
    .X(_18065_));
 sky130_fd_sc_hd__xor2_2 _27884_ (.A(_18059_),
    .B(_18065_),
    .X(_18066_));
 sky130_fd_sc_hd__nand2_2 _27885_ (.A(_18058_),
    .B(_18066_),
    .Y(_18067_));
 sky130_fd_sc_hd__or2_2 _27886_ (.A(_18058_),
    .B(_18066_),
    .X(_18068_));
 sky130_fd_sc_hd__nand2_2 _27887_ (.A(_18067_),
    .B(_18068_),
    .Y(_18069_));
 sky130_fd_sc_hd__a21bo_2 _27888_ (.A1(_17851_),
    .A2(_17857_),
    .B1_N(_17850_),
    .X(_18070_));
 sky130_fd_sc_hd__xnor2_2 _27889_ (.A(_18069_),
    .B(_18070_),
    .Y(_18071_));
 sky130_fd_sc_hd__xnor2_2 _27890_ (.A(_17854_),
    .B(_18071_),
    .Y(_18072_));
 sky130_fd_sc_hd__nand2_2 _27891_ (.A(_17860_),
    .B(_17861_),
    .Y(_18073_));
 sky130_fd_sc_hd__o21a_2 _27892_ (.A1(_17362_),
    .A2(_17862_),
    .B1(_18073_),
    .X(_18074_));
 sky130_fd_sc_hd__xnor2_2 _27893_ (.A(_18072_),
    .B(_18074_),
    .Y(_18076_));
 sky130_fd_sc_hd__xnor2_2 _27894_ (.A(_17948_),
    .B(_18076_),
    .Y(_18077_));
 sky130_fd_sc_hd__nand2_2 _27895_ (.A(_17746_),
    .B(_17864_),
    .Y(_18078_));
 sky130_fd_sc_hd__o21a_2 _27896_ (.A1(_17865_),
    .A2(_17868_),
    .B1(_18078_),
    .X(_18079_));
 sky130_fd_sc_hd__xnor2_2 _27897_ (.A(_18077_),
    .B(_18079_),
    .Y(_18080_));
 sky130_fd_sc_hd__and2b_2 _27898_ (.A_N(_17734_),
    .B(_17733_),
    .X(_18081_));
 sky130_fd_sc_hd__nor2_2 _27899_ (.A(_17610_),
    .B(_17735_),
    .Y(_18082_));
 sky130_fd_sc_hd__or2b_2 _27900_ (.A(_17730_),
    .B_N(_17731_),
    .X(_18083_));
 sky130_fd_sc_hd__or2_4 _27901_ (.A(_17616_),
    .B(_17732_),
    .X(_18084_));
 sky130_fd_sc_hd__and2b_2 _27902_ (.A_N(_17658_),
    .B(_17617_),
    .X(_18085_));
 sky130_fd_sc_hd__a21o_2 _27903_ (.A1(_17619_),
    .A2(_17657_),
    .B1(_18085_),
    .X(_18087_));
 sky130_fd_sc_hd__and2b_2 _27904_ (.A_N(_17640_),
    .B(_17641_),
    .X(_18088_));
 sky130_fd_sc_hd__inv_2 _27905_ (.A(_18088_),
    .Y(_18089_));
 sky130_fd_sc_hd__or2_2 _27906_ (.A(_17634_),
    .B(_17642_),
    .X(_18090_));
 sky130_fd_sc_hd__nor2_2 _27907_ (.A(_17633_),
    .B(_18089_),
    .Y(_18091_));
 sky130_fd_sc_hd__a31o_2 _27908_ (.A1(_17633_),
    .A2(_18089_),
    .A3(_18090_),
    .B1(_18091_),
    .X(_18092_));
 sky130_fd_sc_hd__xnor2_2 _27909_ (.A(_18087_),
    .B(_18092_),
    .Y(_18093_));
 sky130_fd_sc_hd__or2b_2 _27910_ (.A(_17728_),
    .B_N(_17727_),
    .X(_18094_));
 sky130_fd_sc_hd__nand2_2 _27911_ (.A(_17660_),
    .B(_17729_),
    .Y(_18095_));
 sky130_fd_sc_hd__or2_2 _27912_ (.A(_17654_),
    .B(_17655_),
    .X(_18096_));
 sky130_fd_sc_hd__or2_2 _27913_ (.A(_17643_),
    .B(_17656_),
    .X(_18098_));
 sky130_fd_sc_hd__nand2b_2 _27914_ (.A_N(_17680_),
    .B(_17662_),
    .Y(_18099_));
 sky130_fd_sc_hd__or3_2 _27915_ (.A(_12468_),
    .B(_17623_),
    .C(_17625_),
    .X(_18100_));
 sky130_fd_sc_hd__nor2_2 _27916_ (.A(_17623_),
    .B(_17625_),
    .Y(_18101_));
 sky130_fd_sc_hd__a22o_2 _27917_ (.A1(_15616_),
    .A2(_17630_),
    .B1(_18101_),
    .B2(_12838_),
    .X(_18102_));
 sky130_fd_sc_hd__o21a_2 _27918_ (.A1(_17631_),
    .A2(_18100_),
    .B1(_18102_),
    .X(_18103_));
 sky130_fd_sc_hd__inv_2 _27919_ (.A(_17620_),
    .Y(_18104_));
 sky130_fd_sc_hd__or2_2 _27920_ (.A(iY[23]),
    .B(iY[55]),
    .X(_18105_));
 sky130_fd_sc_hd__nand2_2 _27921_ (.A(iY[23]),
    .B(iY[55]),
    .Y(_18106_));
 sky130_fd_sc_hd__nand2_2 _27922_ (.A(_18105_),
    .B(_18106_),
    .Y(_18107_));
 sky130_fd_sc_hd__bufinv_8 _27923_ (.A(_18107_),
    .Y(_18109_));
 sky130_fd_sc_hd__nor3_2 _27924_ (.A(_18104_),
    .B(_17623_),
    .C(_18109_),
    .Y(_18110_));
 sky130_fd_sc_hd__buf_6 _27925_ (.A(_18110_),
    .X(_18111_));
 sky130_fd_sc_hd__o21a_2 _27926_ (.A1(_18104_),
    .A2(_17623_),
    .B1(_18109_),
    .X(_18112_));
 sky130_fd_sc_hd__buf_2 _27927_ (.A(_18112_),
    .X(_18113_));
 sky130_fd_sc_hd__or2_4 _27928_ (.A(_18111_),
    .B(_18113_),
    .X(_18114_));
 sky130_fd_sc_hd__nor2_2 _27929_ (.A(_11578_),
    .B(_18114_),
    .Y(_18115_));
 sky130_fd_sc_hd__xnor2_2 _27930_ (.A(_18103_),
    .B(_18115_),
    .Y(_18116_));
 sky130_fd_sc_hd__o22a_2 _27931_ (.A1(_14640_),
    .A2(_16257_),
    .B1(_16617_),
    .B2(_14346_),
    .X(_18117_));
 sky130_fd_sc_hd__a31o_2 _27932_ (.A1(_15624_),
    .A2(_16613_),
    .A3(_17636_),
    .B1(_18117_),
    .X(_18118_));
 sky130_fd_sc_hd__bufbuf_8 _27933_ (.A(_15167_),
    .X(_18120_));
 sky130_fd_sc_hd__or2_2 _27934_ (.A(_18120_),
    .B(_16922_),
    .X(_18121_));
 sky130_fd_sc_hd__xnor2_2 _27935_ (.A(_18118_),
    .B(_18121_),
    .Y(_18122_));
 sky130_fd_sc_hd__nand2_2 _27936_ (.A(_17635_),
    .B(_17636_),
    .Y(_18123_));
 sky130_fd_sc_hd__o21a_2 _27937_ (.A1(_17638_),
    .A2(_17639_),
    .B1(_18123_),
    .X(_18124_));
 sky130_fd_sc_hd__xnor2_2 _27938_ (.A(_18122_),
    .B(_18124_),
    .Y(_18125_));
 sky130_fd_sc_hd__xor2_2 _27939_ (.A(_18116_),
    .B(_18125_),
    .X(_18126_));
 sky130_fd_sc_hd__nand2_2 _27940_ (.A(_17646_),
    .B(_17652_),
    .Y(_18127_));
 sky130_fd_sc_hd__nand2_2 _27941_ (.A(_17644_),
    .B(_17653_),
    .Y(_18128_));
 sky130_fd_sc_hd__a21bo_2 _27942_ (.A1(_17649_),
    .A2(_17651_),
    .B1_N(_17647_),
    .X(_18129_));
 sky130_fd_sc_hd__a2bb2o_2 _27943_ (.A1_N(_17442_),
    .A2_N(_17664_),
    .B1(_17665_),
    .B2(_17667_),
    .X(_18131_));
 sky130_fd_sc_hd__or4_2 _27944_ (.A(_14357_),
    .B(_14352_),
    .C(_15153_),
    .D(_15597_),
    .X(_18132_));
 sky130_fd_sc_hd__a2bb2o_2 _27945_ (.A1_N(_14357_),
    .A2_N(_15597_),
    .B1(_15585_),
    .B2(_14652_),
    .X(_18133_));
 sky130_fd_sc_hd__nand4_2 _27946_ (.A(_16268_),
    .B(_16933_),
    .C(_18132_),
    .D(_18133_),
    .Y(_18134_));
 sky130_fd_sc_hd__a22o_2 _27947_ (.A1(_16268_),
    .A2(_16933_),
    .B1(_18132_),
    .B2(_18133_),
    .X(_18135_));
 sky130_fd_sc_hd__nand3_2 _27948_ (.A(_18131_),
    .B(_18134_),
    .C(_18135_),
    .Y(_18136_));
 sky130_fd_sc_hd__a21o_2 _27949_ (.A1(_18134_),
    .A2(_18135_),
    .B1(_18131_),
    .X(_18137_));
 sky130_fd_sc_hd__and3_2 _27950_ (.A(_18129_),
    .B(_18136_),
    .C(_18137_),
    .X(_18138_));
 sky130_fd_sc_hd__a21oi_2 _27951_ (.A1(_18136_),
    .A2(_18137_),
    .B1(_18129_),
    .Y(_18139_));
 sky130_fd_sc_hd__or2_2 _27952_ (.A(_18138_),
    .B(_18139_),
    .X(_18140_));
 sky130_fd_sc_hd__a21o_2 _27953_ (.A1(_18127_),
    .A2(_18128_),
    .B1(_18140_),
    .X(_18142_));
 sky130_fd_sc_hd__nand3_2 _27954_ (.A(_18127_),
    .B(_18128_),
    .C(_18140_),
    .Y(_18143_));
 sky130_fd_sc_hd__and3_2 _27955_ (.A(_18126_),
    .B(_18142_),
    .C(_18143_),
    .X(_18144_));
 sky130_fd_sc_hd__a21oi_2 _27956_ (.A1(_18142_),
    .A2(_18143_),
    .B1(_18126_),
    .Y(_18145_));
 sky130_fd_sc_hd__a211oi_2 _27957_ (.A1(_17678_),
    .A2(_18099_),
    .B1(_18144_),
    .C1(_18145_),
    .Y(_18146_));
 sky130_fd_sc_hd__o211a_2 _27958_ (.A1(_18144_),
    .A2(_18145_),
    .B1(_17678_),
    .C1(_18099_),
    .X(_18147_));
 sky130_fd_sc_hd__a211oi_2 _27959_ (.A1(_18096_),
    .A2(_18098_),
    .B1(_18146_),
    .C1(_18147_),
    .Y(_18148_));
 sky130_fd_sc_hd__o211a_2 _27960_ (.A1(_18146_),
    .A2(_18147_),
    .B1(_18096_),
    .C1(_18098_),
    .X(_18149_));
 sky130_fd_sc_hd__or2b_2 _27961_ (.A(_17723_),
    .B_N(_17724_),
    .X(_18150_));
 sky130_fd_sc_hd__nand2_2 _27962_ (.A(_17682_),
    .B(_17726_),
    .Y(_18151_));
 sky130_fd_sc_hd__or2_2 _27963_ (.A(_17673_),
    .B(_17675_),
    .X(_18153_));
 sky130_fd_sc_hd__o21ai_2 _27964_ (.A1(_17668_),
    .A2(_17676_),
    .B1(_18153_),
    .Y(_18154_));
 sky130_fd_sc_hd__a21oi_2 _27965_ (.A1(_17683_),
    .A2(_17693_),
    .B1(_17691_),
    .Y(_18155_));
 sky130_fd_sc_hd__or4_2 _27966_ (.A(_15211_),
    .B(_15647_),
    .C(_15168_),
    .D(_15169_),
    .X(_18156_));
 sky130_fd_sc_hd__buf_1 _27967_ (.A(_13938_),
    .X(_18157_));
 sky130_fd_sc_hd__a22o_2 _27968_ (.A1(_18157_),
    .A2(_14410_),
    .B1(_14605_),
    .B2(_13845_),
    .X(_18158_));
 sky130_fd_sc_hd__nor2_2 _27969_ (.A(_14983_),
    .B(_14948_),
    .Y(_18159_));
 sky130_fd_sc_hd__and3_2 _27970_ (.A(_18156_),
    .B(_18158_),
    .C(_18159_),
    .X(_18160_));
 sky130_fd_sc_hd__a21oi_2 _27971_ (.A1(_18156_),
    .A2(_18158_),
    .B1(_18159_),
    .Y(_18161_));
 sky130_fd_sc_hd__or2_2 _27972_ (.A(_18160_),
    .B(_18161_),
    .X(_18162_));
 sky130_fd_sc_hd__and3_2 _27973_ (.A(_13887_),
    .B(_14995_),
    .C(_14996_),
    .X(_18164_));
 sky130_fd_sc_hd__a32o_2 _27974_ (.A1(_13542_),
    .A2(_14995_),
    .A3(_14996_),
    .B1(_13888_),
    .B2(_14999_),
    .X(_18165_));
 sky130_fd_sc_hd__a21bo_2 _27975_ (.A1(_17669_),
    .A2(_18164_),
    .B1_N(_18165_),
    .X(_18166_));
 sky130_fd_sc_hd__nor2_2 _27976_ (.A(_13972_),
    .B(_14988_),
    .Y(_18167_));
 sky130_fd_sc_hd__xor2_2 _27977_ (.A(_18166_),
    .B(_18167_),
    .X(_18168_));
 sky130_fd_sc_hd__o2bb2a_2 _27978_ (.A1_N(_17446_),
    .A2_N(_17669_),
    .B1(_17671_),
    .B2(_17672_),
    .X(_18169_));
 sky130_fd_sc_hd__xnor2_2 _27979_ (.A(_18168_),
    .B(_18169_),
    .Y(_18170_));
 sky130_fd_sc_hd__xnor2_2 _27980_ (.A(_18162_),
    .B(_18170_),
    .Y(_18171_));
 sky130_fd_sc_hd__xnor2_2 _27981_ (.A(_18155_),
    .B(_18171_),
    .Y(_18172_));
 sky130_fd_sc_hd__xnor2_2 _27982_ (.A(_18154_),
    .B(_18172_),
    .Y(_18173_));
 sky130_fd_sc_hd__or2_2 _27983_ (.A(_17720_),
    .B(_17721_),
    .X(_18175_));
 sky130_fd_sc_hd__nand2_2 _27984_ (.A(_17695_),
    .B(_17722_),
    .Y(_18176_));
 sky130_fd_sc_hd__nand2_2 _27985_ (.A(_17687_),
    .B(_17689_),
    .Y(_18177_));
 sky130_fd_sc_hd__or4_4 _27986_ (.A(_15650_),
    .B(_14978_),
    .C(_16988_),
    .D(_17007_),
    .X(_18178_));
 sky130_fd_sc_hd__o31a_2 _27987_ (.A1(_14356_),
    .A2(_17696_),
    .A3(_17699_),
    .B1(_18178_),
    .X(_18179_));
 sky130_fd_sc_hd__nand2_2 _27988_ (.A(_15223_),
    .B(_15225_),
    .Y(_18180_));
 sky130_fd_sc_hd__buf_1 _27989_ (.A(_18180_),
    .X(_18181_));
 sky130_fd_sc_hd__nor2_2 _27990_ (.A(_12773_),
    .B(_16677_),
    .Y(_18182_));
 sky130_fd_sc_hd__xnor2_2 _27991_ (.A(_17686_),
    .B(_18182_),
    .Y(_18183_));
 sky130_fd_sc_hd__nor3_2 _27992_ (.A(_14625_),
    .B(_18181_),
    .C(_18183_),
    .Y(_18184_));
 sky130_fd_sc_hd__o21a_2 _27993_ (.A1(_14625_),
    .A2(_18181_),
    .B1(_18183_),
    .X(_18186_));
 sky130_fd_sc_hd__or3_4 _27994_ (.A(_18179_),
    .B(_18184_),
    .C(_18186_),
    .X(_18187_));
 sky130_fd_sc_hd__o21ai_2 _27995_ (.A1(_18184_),
    .A2(_18186_),
    .B1(_18179_),
    .Y(_18188_));
 sky130_fd_sc_hd__and3_2 _27996_ (.A(_18177_),
    .B(_18187_),
    .C(_18188_),
    .X(_18189_));
 sky130_fd_sc_hd__a21oi_2 _27997_ (.A1(_18187_),
    .A2(_18188_),
    .B1(_18177_),
    .Y(_18190_));
 sky130_fd_sc_hd__or2_4 _27998_ (.A(_18189_),
    .B(_18190_),
    .X(_18191_));
 sky130_fd_sc_hd__buf_1 _27999_ (.A(_12759_),
    .X(_18192_));
 sky130_fd_sc_hd__nand2_2 _28000_ (.A(_18192_),
    .B(_17006_),
    .Y(_18193_));
 sky130_fd_sc_hd__nor2_2 _28001_ (.A(_13926_),
    .B(_16999_),
    .Y(_18194_));
 sky130_fd_sc_hd__and3_2 _28002_ (.A(_14980_),
    .B(_17488_),
    .C(_18194_),
    .X(_18195_));
 sky130_fd_sc_hd__a21o_2 _28003_ (.A1(_14980_),
    .A2(_17488_),
    .B1(_18194_),
    .X(_18197_));
 sky130_fd_sc_hd__and2b_2 _28004_ (.A_N(_18195_),
    .B(_18197_),
    .X(_18198_));
 sky130_fd_sc_hd__xnor2_2 _28005_ (.A(_18193_),
    .B(_18198_),
    .Y(_18199_));
 sky130_fd_sc_hd__buf_1 _28006_ (.A(_17482_),
    .X(_18200_));
 sky130_fd_sc_hd__xnor2_2 _28007_ (.A(iX[23]),
    .B(iX[55]),
    .Y(_18201_));
 sky130_fd_sc_hd__a21oi_4 _28008_ (.A1(_17707_),
    .A2(_17711_),
    .B1(_17708_),
    .Y(_18202_));
 sky130_fd_sc_hd__xor2_2 _28009_ (.A(_18201_),
    .B(_18202_),
    .X(_18203_));
 sky130_fd_sc_hd__and3_4 _28010_ (.A(_11585_),
    .B(_17715_),
    .C(_18203_),
    .X(_18204_));
 sky130_fd_sc_hd__and2_2 _28011_ (.A(_17712_),
    .B(_17713_),
    .X(_18205_));
 sky130_fd_sc_hd__a22o_4 _28012_ (.A1(_11585_),
    .A2(_18205_),
    .B1(_18203_),
    .B2(_11381_),
    .X(_18206_));
 sky130_fd_sc_hd__or4b_4 _28013_ (.A(_11793_),
    .B(_18200_),
    .C(_18204_),
    .D_N(_18206_),
    .X(_18208_));
 sky130_fd_sc_hd__buf_4 _28014_ (.A(_17485_),
    .X(_18209_));
 sky130_fd_sc_hd__xnor2_2 _28015_ (.A(_18201_),
    .B(_18202_),
    .Y(_18210_));
 sky130_fd_sc_hd__buf_2 _28016_ (.A(_18210_),
    .X(_18211_));
 sky130_fd_sc_hd__or3b_4 _28017_ (.A(_11576_),
    .B(_18211_),
    .C_N(_17715_),
    .X(_18212_));
 sky130_fd_sc_hd__a22o_2 _28018_ (.A1(_15677_),
    .A2(_18209_),
    .B1(_18212_),
    .B2(_18206_),
    .X(_18213_));
 sky130_fd_sc_hd__and3_2 _28019_ (.A(_11585_),
    .B(_18209_),
    .C(_17715_),
    .X(_18214_));
 sky130_fd_sc_hd__a31o_2 _28020_ (.A1(_15677_),
    .A2(_17702_),
    .A3(_17716_),
    .B1(_18214_),
    .X(_18215_));
 sky130_fd_sc_hd__nand3_2 _28021_ (.A(_18208_),
    .B(_18213_),
    .C(_18215_),
    .Y(_18216_));
 sky130_fd_sc_hd__a21o_2 _28022_ (.A1(_18208_),
    .A2(_18213_),
    .B1(_18215_),
    .X(_18217_));
 sky130_fd_sc_hd__nand3_2 _28023_ (.A(_18199_),
    .B(_18216_),
    .C(_18217_),
    .Y(_18219_));
 sky130_fd_sc_hd__a21o_2 _28024_ (.A1(_18216_),
    .A2(_18217_),
    .B1(_18199_),
    .X(_18220_));
 sky130_fd_sc_hd__and2b_2 _28025_ (.A_N(_17718_),
    .B(_17717_),
    .X(_18221_));
 sky130_fd_sc_hd__a21o_2 _28026_ (.A1(_17701_),
    .A2(_17719_),
    .B1(_18221_),
    .X(_18222_));
 sky130_fd_sc_hd__and3_2 _28027_ (.A(_18219_),
    .B(_18220_),
    .C(_18222_),
    .X(_18223_));
 sky130_fd_sc_hd__a21oi_2 _28028_ (.A1(_18219_),
    .A2(_18220_),
    .B1(_18222_),
    .Y(_18224_));
 sky130_fd_sc_hd__nor3_2 _28029_ (.A(_18191_),
    .B(_18223_),
    .C(_18224_),
    .Y(_18225_));
 sky130_fd_sc_hd__o21a_2 _28030_ (.A1(_18223_),
    .A2(_18224_),
    .B1(_18191_),
    .X(_18226_));
 sky130_fd_sc_hd__a211o_2 _28031_ (.A1(_18175_),
    .A2(_18176_),
    .B1(_18225_),
    .C1(_18226_),
    .X(_18227_));
 sky130_fd_sc_hd__o211ai_2 _28032_ (.A1(_18225_),
    .A2(_18226_),
    .B1(_18175_),
    .C1(_18176_),
    .Y(_18228_));
 sky130_fd_sc_hd__and3_4 _28033_ (.A(_18173_),
    .B(_18227_),
    .C(_18228_),
    .X(_18230_));
 sky130_fd_sc_hd__a21oi_2 _28034_ (.A1(_18227_),
    .A2(_18228_),
    .B1(_18173_),
    .Y(_18231_));
 sky130_fd_sc_hd__a211oi_4 _28035_ (.A1(_18150_),
    .A2(_18151_),
    .B1(_18230_),
    .C1(_18231_),
    .Y(_18232_));
 sky130_fd_sc_hd__o211a_2 _28036_ (.A1(_18230_),
    .A2(_18231_),
    .B1(_18150_),
    .C1(_18151_),
    .X(_18233_));
 sky130_fd_sc_hd__nor4_2 _28037_ (.A(_18148_),
    .B(_18149_),
    .C(_18232_),
    .D(_18233_),
    .Y(_18234_));
 sky130_fd_sc_hd__o22a_2 _28038_ (.A1(_18148_),
    .A2(_18149_),
    .B1(_18232_),
    .B2(_18233_),
    .X(_18235_));
 sky130_fd_sc_hd__a211o_2 _28039_ (.A1(_18094_),
    .A2(_18095_),
    .B1(_18234_),
    .C1(_18235_),
    .X(_18236_));
 sky130_fd_sc_hd__o211ai_2 _28040_ (.A1(_18234_),
    .A2(_18235_),
    .B1(_18094_),
    .C1(_18095_),
    .Y(_18237_));
 sky130_fd_sc_hd__and3_4 _28041_ (.A(_18093_),
    .B(_18236_),
    .C(_18237_),
    .X(_18238_));
 sky130_fd_sc_hd__a21oi_2 _28042_ (.A1(_18236_),
    .A2(_18237_),
    .B1(_18093_),
    .Y(_18239_));
 sky130_fd_sc_hd__a211o_2 _28043_ (.A1(_18083_),
    .A2(_18084_),
    .B1(_18238_),
    .C1(_18239_),
    .X(_18241_));
 sky130_fd_sc_hd__o211ai_2 _28044_ (.A1(_18238_),
    .A2(_18239_),
    .B1(_18083_),
    .C1(_18084_),
    .Y(_18242_));
 sky130_fd_sc_hd__nand3_2 _28045_ (.A(_17613_),
    .B(_18241_),
    .C(_18242_),
    .Y(_18243_));
 sky130_fd_sc_hd__a21o_2 _28046_ (.A1(_18241_),
    .A2(_18242_),
    .B1(_17613_),
    .X(_18244_));
 sky130_fd_sc_hd__o211ai_2 _28047_ (.A1(_18081_),
    .A2(_18082_),
    .B1(_18243_),
    .C1(_18244_),
    .Y(_18245_));
 sky130_fd_sc_hd__a211o_2 _28048_ (.A1(_18243_),
    .A2(_18244_),
    .B1(_18081_),
    .C1(_18082_),
    .X(_18246_));
 sky130_fd_sc_hd__and2_2 _28049_ (.A(_17609_),
    .B(_17737_),
    .X(_18247_));
 sky130_fd_sc_hd__a21o_2 _28050_ (.A1(_18245_),
    .A2(_18246_),
    .B1(_18247_),
    .X(_18248_));
 sky130_fd_sc_hd__nand2_2 _28051_ (.A(_17609_),
    .B(_17737_),
    .Y(_18249_));
 sky130_fd_sc_hd__nand2_2 _28052_ (.A(_18245_),
    .B(_18246_),
    .Y(_18250_));
 sky130_fd_sc_hd__or2_2 _28053_ (.A(_18249_),
    .B(_18250_),
    .X(_18252_));
 sky130_fd_sc_hd__nand2_2 _28054_ (.A(_18248_),
    .B(_18252_),
    .Y(_18253_));
 sky130_fd_sc_hd__nand2_2 _28055_ (.A(_17608_),
    .B(_17738_),
    .Y(_18254_));
 sky130_fd_sc_hd__a21boi_2 _28056_ (.A1(_17740_),
    .A2(_17743_),
    .B1_N(_18254_),
    .Y(_18255_));
 sky130_fd_sc_hd__xnor2_2 _28057_ (.A(_18253_),
    .B(_18255_),
    .Y(_18256_));
 sky130_fd_sc_hd__xnor2_2 _28058_ (.A(_18080_),
    .B(_18256_),
    .Y(_18257_));
 sky130_fd_sc_hd__xnor2_2 _28059_ (.A(_08066_),
    .B(_18257_),
    .Y(_18258_));
 sky130_fd_sc_hd__and3_2 _28060_ (.A(_17946_),
    .B(_17947_),
    .C(_18258_),
    .X(_18259_));
 sky130_fd_sc_hd__a21oi_2 _28061_ (.A1(_17946_),
    .A2(_17947_),
    .B1(_18258_),
    .Y(_18260_));
 sky130_fd_sc_hd__nor2_2 _28062_ (.A(_18259_),
    .B(_18260_),
    .Y(_18261_));
 sky130_fd_sc_hd__xnor2_2 _28063_ (.A(_17945_),
    .B(_18261_),
    .Y(_18263_));
 sky130_fd_sc_hd__xor2_2 _28064_ (.A(_17944_),
    .B(_18263_),
    .X(_18264_));
 sky130_fd_sc_hd__o21ba_2 _28065_ (.A1(_17884_),
    .A2(_17888_),
    .B1_N(_17883_),
    .X(_18265_));
 sky130_fd_sc_hd__xnor2_2 _28066_ (.A(_18264_),
    .B(_18265_),
    .Y(oO[55]));
 sky130_fd_sc_hd__nor2_2 _28067_ (.A(_17602_),
    .B(_17941_),
    .Y(_18266_));
 sky130_fd_sc_hd__or2_2 _28068_ (.A(_17191_),
    .B(_17256_),
    .X(_18267_));
 sky130_fd_sc_hd__and3b_2 _28069_ (.A_N(_17257_),
    .B(_18266_),
    .C(_18267_),
    .X(_18268_));
 sky130_fd_sc_hd__a21oi_2 _28070_ (.A1(_17600_),
    .A2(_17940_),
    .B1(_17939_),
    .Y(_18269_));
 sky130_fd_sc_hd__a311o_2 _28071_ (.A1(_16888_),
    .A2(_17258_),
    .A3(_18266_),
    .B1(_18268_),
    .C1(_18269_),
    .X(_18270_));
 sky130_fd_sc_hd__nand2_2 _28072_ (.A(_17930_),
    .B(_17931_),
    .Y(_18271_));
 sky130_fd_sc_hd__or2b_2 _28073_ (.A(_17914_),
    .B_N(_17913_),
    .X(_18273_));
 sky130_fd_sc_hd__and4_2 _28074_ (.A(iY[27]),
    .B(iX[28]),
    .C(iY[28]),
    .D(iX[29]),
    .X(_18274_));
 sky130_fd_sc_hd__a22oi_2 _28075_ (.A1(iX[28]),
    .A2(iY[28]),
    .B1(iX[29]),
    .B2(iY[27]),
    .Y(_18275_));
 sky130_fd_sc_hd__nor2_2 _28076_ (.A(_18274_),
    .B(_18275_),
    .Y(_18276_));
 sky130_fd_sc_hd__nand2_2 _28077_ (.A(iX[27]),
    .B(iY[29]),
    .Y(_18277_));
 sky130_fd_sc_hd__xnor2_2 _28078_ (.A(_18276_),
    .B(_18277_),
    .Y(_18278_));
 sky130_fd_sc_hd__o21ba_2 _28079_ (.A1(_17909_),
    .A2(_17912_),
    .B1_N(_17908_),
    .X(_18279_));
 sky130_fd_sc_hd__xnor2_2 _28080_ (.A(_18278_),
    .B(_18279_),
    .Y(_18280_));
 sky130_fd_sc_hd__nand3_2 _28081_ (.A(iX[26]),
    .B(iY[30]),
    .C(_18280_),
    .Y(_18281_));
 sky130_fd_sc_hd__a21o_2 _28082_ (.A1(iX[26]),
    .A2(iY[30]),
    .B1(_18280_),
    .X(_18282_));
 sky130_fd_sc_hd__nand2_2 _28083_ (.A(_18281_),
    .B(_18282_),
    .Y(_18284_));
 sky130_fd_sc_hd__a21o_2 _28084_ (.A1(_18273_),
    .A2(_17916_),
    .B1(_18284_),
    .X(_18285_));
 sky130_fd_sc_hd__nand3_2 _28085_ (.A(_18273_),
    .B(_17916_),
    .C(_18284_),
    .Y(_18286_));
 sky130_fd_sc_hd__and2_2 _28086_ (.A(_18285_),
    .B(_18286_),
    .X(_18287_));
 sky130_fd_sc_hd__a21o_2 _28087_ (.A1(iX[25]),
    .A2(iY[31]),
    .B1(_18287_),
    .X(_18288_));
 sky130_fd_sc_hd__nand3_2 _28088_ (.A(iX[25]),
    .B(iY[31]),
    .C(_18287_),
    .Y(_18289_));
 sky130_fd_sc_hd__and2_2 _28089_ (.A(_18288_),
    .B(_18289_),
    .X(_18290_));
 sky130_fd_sc_hd__a31o_2 _28090_ (.A1(iY[26]),
    .A2(iX[29]),
    .A3(_17892_),
    .B1(_17891_),
    .X(_18291_));
 sky130_fd_sc_hd__a22oi_2 _28091_ (.A1(iY[26]),
    .A2(iX[30]),
    .B1(iX[31]),
    .B2(iY[25]),
    .Y(_18292_));
 sky130_fd_sc_hd__and4_2 _28092_ (.A(iY[25]),
    .B(iY[26]),
    .C(iX[30]),
    .D(iX[31]),
    .X(_18293_));
 sky130_fd_sc_hd__nor2_2 _28093_ (.A(_18292_),
    .B(_18293_),
    .Y(_18295_));
 sky130_fd_sc_hd__and2_2 _28094_ (.A(_18291_),
    .B(_18295_),
    .X(_18296_));
 sky130_fd_sc_hd__nor2_2 _28095_ (.A(_18291_),
    .B(_18295_),
    .Y(_18297_));
 sky130_fd_sc_hd__nor2_2 _28096_ (.A(_18296_),
    .B(_18297_),
    .Y(_18298_));
 sky130_fd_sc_hd__a21oi_2 _28097_ (.A1(_17896_),
    .A2(_17897_),
    .B1(_17901_),
    .Y(_18299_));
 sky130_fd_sc_hd__xnor2_2 _28098_ (.A(_18298_),
    .B(_18299_),
    .Y(_18300_));
 sky130_fd_sc_hd__xnor2_2 _28099_ (.A(_18290_),
    .B(_18300_),
    .Y(_18301_));
 sky130_fd_sc_hd__a21oi_2 _28100_ (.A1(_17905_),
    .A2(_17926_),
    .B1(_18301_),
    .Y(_18302_));
 sky130_fd_sc_hd__nand3_2 _28101_ (.A(_17905_),
    .B(_17926_),
    .C(_18301_),
    .Y(_18303_));
 sky130_fd_sc_hd__or2b_2 _28102_ (.A(_18302_),
    .B_N(_18303_),
    .X(_18304_));
 sky130_fd_sc_hd__xnor2_2 _28103_ (.A(_17928_),
    .B(_18304_),
    .Y(_18306_));
 sky130_fd_sc_hd__xnor2_2 _28104_ (.A(_18271_),
    .B(_18306_),
    .Y(_18307_));
 sky130_fd_sc_hd__a31o_2 _28105_ (.A1(iX[24]),
    .A2(iY[31]),
    .A3(_17922_),
    .B1(_17919_),
    .X(_18308_));
 sky130_fd_sc_hd__xnor2_2 _28106_ (.A(_18307_),
    .B(_18308_),
    .Y(_18309_));
 sky130_fd_sc_hd__a21o_2 _28107_ (.A1(_17890_),
    .A2(_17933_),
    .B1(_17936_),
    .X(_18310_));
 sky130_fd_sc_hd__xnor2_2 _28108_ (.A(_18309_),
    .B(_18310_),
    .Y(_18311_));
 sky130_fd_sc_hd__xnor2_2 _28109_ (.A(_18270_),
    .B(_18311_),
    .Y(_18312_));
 sky130_fd_sc_hd__and3_2 _28110_ (.A(_18247_),
    .B(_18245_),
    .C(_18246_),
    .X(_18313_));
 sky130_fd_sc_hd__or3b_4 _28111_ (.A(_18313_),
    .B(_17739_),
    .C_N(_18248_),
    .X(_18314_));
 sky130_fd_sc_hd__or2b_2 _28112_ (.A(_18314_),
    .B_N(_17742_),
    .X(_18315_));
 sky130_fd_sc_hd__a21o_2 _28113_ (.A1(_18249_),
    .A2(_18254_),
    .B1(_18250_),
    .X(_18317_));
 sky130_fd_sc_hd__o41a_2 _28114_ (.A1(_17521_),
    .A2(_17522_),
    .A3(_17519_),
    .A4(_18314_),
    .B1(_18317_),
    .X(_18318_));
 sky130_fd_sc_hd__nand2_2 _28115_ (.A(_18315_),
    .B(_18318_),
    .Y(_18319_));
 sky130_fd_sc_hd__inv_2 _28116_ (.A(_18241_),
    .Y(_18320_));
 sky130_fd_sc_hd__and3_2 _28117_ (.A(_17613_),
    .B(_18241_),
    .C(_18242_),
    .X(_18321_));
 sky130_fd_sc_hd__and2b_2 _28118_ (.A_N(_18092_),
    .B(_18087_),
    .X(_18322_));
 sky130_fd_sc_hd__inv_2 _28119_ (.A(_18236_),
    .Y(_18323_));
 sky130_fd_sc_hd__or2_2 _28120_ (.A(_18122_),
    .B(_18124_),
    .X(_18324_));
 sky130_fd_sc_hd__o21ai_2 _28121_ (.A1(_18116_),
    .A2(_18125_),
    .B1(_18324_),
    .Y(_18325_));
 sky130_fd_sc_hd__nor2_2 _28122_ (.A(_18111_),
    .B(_18113_),
    .Y(_18326_));
 sky130_fd_sc_hd__buf_2 _28123_ (.A(_18326_),
    .X(_18328_));
 sky130_fd_sc_hd__nor2_2 _28124_ (.A(_17631_),
    .B(_18100_),
    .Y(_18329_));
 sky130_fd_sc_hd__a31o_2 _28125_ (.A1(_14592_),
    .A2(_18102_),
    .A3(_18328_),
    .B1(_18329_),
    .X(_18330_));
 sky130_fd_sc_hd__nand2_2 _28126_ (.A(iY[24]),
    .B(iY[56]),
    .Y(_18331_));
 sky130_fd_sc_hd__or2_2 _28127_ (.A(iY[24]),
    .B(iY[56]),
    .X(_18332_));
 sky130_fd_sc_hd__nand2_2 _28128_ (.A(_18331_),
    .B(_18332_),
    .Y(_18333_));
 sky130_fd_sc_hd__or2_2 _28129_ (.A(_17622_),
    .B(_18107_),
    .X(_18334_));
 sky130_fd_sc_hd__nand2_2 _28130_ (.A(_17620_),
    .B(_18106_),
    .Y(_18335_));
 sky130_fd_sc_hd__o2bb2a_2 _28131_ (.A1_N(_18105_),
    .A2_N(_18335_),
    .B1(_18334_),
    .B2(_17624_),
    .X(_18336_));
 sky130_fd_sc_hd__o31a_2 _28132_ (.A1(_16920_),
    .A2(_17403_),
    .A3(_18334_),
    .B1(_18336_),
    .X(_18337_));
 sky130_fd_sc_hd__and3_4 _28133_ (.A(_16912_),
    .B(_16916_),
    .C(_18336_),
    .X(_18339_));
 sky130_fd_sc_hd__or3_4 _28134_ (.A(_18333_),
    .B(_18337_),
    .C(_18339_),
    .X(_18340_));
 sky130_fd_sc_hd__o21ai_2 _28135_ (.A1(_18337_),
    .A2(_18339_),
    .B1(_18333_),
    .Y(_18341_));
 sky130_fd_sc_hd__nand2_2 _28136_ (.A(_18340_),
    .B(_18341_),
    .Y(_18342_));
 sky130_fd_sc_hd__buf_2 _28137_ (.A(_18342_),
    .X(_18343_));
 sky130_fd_sc_hd__buf_1 _28138_ (.A(_18343_),
    .X(_18344_));
 sky130_fd_sc_hd__nor2_2 _28139_ (.A(_11579_),
    .B(_18344_),
    .Y(_18345_));
 sky130_fd_sc_hd__xnor2_2 _28140_ (.A(_18330_),
    .B(_18345_),
    .Y(_18346_));
 sky130_fd_sc_hd__xnor2_2 _28141_ (.A(_18325_),
    .B(_18346_),
    .Y(_18347_));
 sky130_fd_sc_hd__and2_2 _28142_ (.A(_18091_),
    .B(_18347_),
    .X(_18348_));
 sky130_fd_sc_hd__nor2_2 _28143_ (.A(_18091_),
    .B(_18347_),
    .Y(_18350_));
 sky130_fd_sc_hd__nor2_2 _28144_ (.A(_18348_),
    .B(_18350_),
    .Y(_18351_));
 sky130_fd_sc_hd__o21ai_2 _28145_ (.A1(_18146_),
    .A2(_18148_),
    .B1(_18351_),
    .Y(_18352_));
 sky130_fd_sc_hd__or3_2 _28146_ (.A(_18146_),
    .B(_18148_),
    .C(_18351_),
    .X(_18353_));
 sky130_fd_sc_hd__and2_2 _28147_ (.A(_18352_),
    .B(_18353_),
    .X(_18354_));
 sky130_fd_sc_hd__a21bo_2 _28148_ (.A1(_18126_),
    .A2(_18143_),
    .B1_N(_18142_),
    .X(_18355_));
 sky130_fd_sc_hd__nor2_2 _28149_ (.A(_18155_),
    .B(_18171_),
    .Y(_18356_));
 sky130_fd_sc_hd__and2b_2 _28150_ (.A_N(_18172_),
    .B(_18154_),
    .X(_18357_));
 sky130_fd_sc_hd__or3_4 _28151_ (.A(_15167_),
    .B(_17404_),
    .C(_17405_),
    .X(_18358_));
 sky130_fd_sc_hd__xor2_2 _28152_ (.A(_18100_),
    .B(_18358_),
    .X(_18359_));
 sky130_fd_sc_hd__or3_2 _28153_ (.A(_11571_),
    .B(_18111_),
    .C(_18113_),
    .X(_18361_));
 sky130_fd_sc_hd__xnor2_2 _28154_ (.A(_18359_),
    .B(_18361_),
    .Y(_18362_));
 sky130_fd_sc_hd__buf_1 _28155_ (.A(_16922_),
    .X(_18363_));
 sky130_fd_sc_hd__nor2_2 _28156_ (.A(_14343_),
    .B(_16255_),
    .Y(_18364_));
 sky130_fd_sc_hd__and3_2 _28157_ (.A(_15624_),
    .B(_16613_),
    .C(_18364_),
    .X(_18365_));
 sky130_fd_sc_hd__a21o_2 _28158_ (.A1(_15624_),
    .A2(_16613_),
    .B1(_18364_),
    .X(_18366_));
 sky130_fd_sc_hd__or4b_2 _28159_ (.A(_16271_),
    .B(_18363_),
    .C(_18365_),
    .D_N(_18366_),
    .X(_18367_));
 sky130_fd_sc_hd__buf_1 _28160_ (.A(_14640_),
    .X(_18368_));
 sky130_fd_sc_hd__or3b_2 _28161_ (.A(_18368_),
    .B(_16617_),
    .C_N(_18364_),
    .X(_18369_));
 sky130_fd_sc_hd__a22o_2 _28162_ (.A1(_14629_),
    .A2(_17394_),
    .B1(_18369_),
    .B2(_18366_),
    .X(_18370_));
 sky130_fd_sc_hd__or3b_2 _28163_ (.A(_18368_),
    .B(_16619_),
    .C_N(_17636_),
    .X(_18372_));
 sky130_fd_sc_hd__o21ai_2 _28164_ (.A1(_18117_),
    .A2(_18121_),
    .B1(_18372_),
    .Y(_18373_));
 sky130_fd_sc_hd__nand3_2 _28165_ (.A(_18367_),
    .B(_18370_),
    .C(_18373_),
    .Y(_18374_));
 sky130_fd_sc_hd__a21o_2 _28166_ (.A1(_18367_),
    .A2(_18370_),
    .B1(_18373_),
    .X(_18375_));
 sky130_fd_sc_hd__nand3_2 _28167_ (.A(_18362_),
    .B(_18374_),
    .C(_18375_),
    .Y(_18376_));
 sky130_fd_sc_hd__a21o_2 _28168_ (.A1(_18374_),
    .A2(_18375_),
    .B1(_18362_),
    .X(_18377_));
 sky130_fd_sc_hd__nand2_2 _28169_ (.A(_18132_),
    .B(_18134_),
    .Y(_18378_));
 sky130_fd_sc_hd__a21bo_2 _28170_ (.A1(_18158_),
    .A2(_18159_),
    .B1_N(_18156_),
    .X(_18379_));
 sky130_fd_sc_hd__or2_2 _28171_ (.A(_14983_),
    .B(_15596_),
    .X(_18380_));
 sky130_fd_sc_hd__or3_2 _28172_ (.A(_14352_),
    .B(_16237_),
    .C(_18380_),
    .X(_18381_));
 sky130_fd_sc_hd__a2bb2o_2 _28173_ (.A1_N(_14352_),
    .A2_N(_15598_),
    .B1(_15586_),
    .B2(_14648_),
    .X(_18383_));
 sky130_fd_sc_hd__nor2_2 _28174_ (.A(_14357_),
    .B(_15834_),
    .Y(_18384_));
 sky130_fd_sc_hd__nand3_2 _28175_ (.A(_18381_),
    .B(_18383_),
    .C(_18384_),
    .Y(_18385_));
 sky130_fd_sc_hd__a21o_2 _28176_ (.A1(_18381_),
    .A2(_18383_),
    .B1(_18384_),
    .X(_18386_));
 sky130_fd_sc_hd__nand3_2 _28177_ (.A(_18379_),
    .B(_18385_),
    .C(_18386_),
    .Y(_18387_));
 sky130_fd_sc_hd__a21o_2 _28178_ (.A1(_18385_),
    .A2(_18386_),
    .B1(_18379_),
    .X(_18388_));
 sky130_fd_sc_hd__nand3_2 _28179_ (.A(_18378_),
    .B(_18387_),
    .C(_18388_),
    .Y(_18389_));
 sky130_fd_sc_hd__a21o_2 _28180_ (.A1(_18387_),
    .A2(_18388_),
    .B1(_18378_),
    .X(_18390_));
 sky130_fd_sc_hd__a21bo_2 _28181_ (.A1(_18129_),
    .A2(_18137_),
    .B1_N(_18136_),
    .X(_18391_));
 sky130_fd_sc_hd__nand3_2 _28182_ (.A(_18389_),
    .B(_18390_),
    .C(_18391_),
    .Y(_18392_));
 sky130_fd_sc_hd__a21o_2 _28183_ (.A1(_18389_),
    .A2(_18390_),
    .B1(_18391_),
    .X(_18394_));
 sky130_fd_sc_hd__nand4_2 _28184_ (.A(_18376_),
    .B(_18377_),
    .C(_18392_),
    .D(_18394_),
    .Y(_18395_));
 sky130_fd_sc_hd__a22o_2 _28185_ (.A1(_18376_),
    .A2(_18377_),
    .B1(_18392_),
    .B2(_18394_),
    .X(_18396_));
 sky130_fd_sc_hd__o211a_2 _28186_ (.A1(_18356_),
    .A2(_18357_),
    .B1(_18395_),
    .C1(_18396_),
    .X(_18397_));
 sky130_fd_sc_hd__a211oi_2 _28187_ (.A1(_18395_),
    .A2(_18396_),
    .B1(_18356_),
    .C1(_18357_),
    .Y(_18398_));
 sky130_fd_sc_hd__nor2_2 _28188_ (.A(_18397_),
    .B(_18398_),
    .Y(_18399_));
 sky130_fd_sc_hd__xor2_2 _28189_ (.A(_18355_),
    .B(_18399_),
    .X(_18400_));
 sky130_fd_sc_hd__nand3_2 _28190_ (.A(_18173_),
    .B(_18227_),
    .C(_18228_),
    .Y(_18401_));
 sky130_fd_sc_hd__o32a_2 _28191_ (.A1(_18160_),
    .A2(_18161_),
    .A3(_18170_),
    .B1(_18169_),
    .B2(_18168_),
    .X(_18402_));
 sky130_fd_sc_hd__a21bo_2 _28192_ (.A1(_18177_),
    .A2(_18188_),
    .B1_N(_18187_),
    .X(_18403_));
 sky130_fd_sc_hd__nand2_2 _28193_ (.A(_15208_),
    .B(_14409_),
    .Y(_18405_));
 sky130_fd_sc_hd__or3_2 _28194_ (.A(_15647_),
    .B(_15169_),
    .C(_18405_),
    .X(_18406_));
 sky130_fd_sc_hd__o21ai_2 _28195_ (.A1(_15647_),
    .A2(_15169_),
    .B1(_18405_),
    .Y(_18407_));
 sky130_fd_sc_hd__and2_2 _28196_ (.A(_18406_),
    .B(_18407_),
    .X(_18408_));
 sky130_fd_sc_hd__nor2_2 _28197_ (.A(_15211_),
    .B(_15173_),
    .Y(_18409_));
 sky130_fd_sc_hd__xnor2_2 _28198_ (.A(_18408_),
    .B(_18409_),
    .Y(_18410_));
 sky130_fd_sc_hd__nor2_2 _28199_ (.A(_13972_),
    .B(_15005_),
    .Y(_18411_));
 sky130_fd_sc_hd__or4b_4 _28200_ (.A(_14612_),
    .B(_15219_),
    .C(_15220_),
    .D_N(_18164_),
    .X(_18412_));
 sky130_fd_sc_hd__a31o_2 _28201_ (.A1(_13543_),
    .A2(_15224_),
    .A3(_15226_),
    .B1(_18164_),
    .X(_18413_));
 sky130_fd_sc_hd__nand3_2 _28202_ (.A(_18411_),
    .B(_18412_),
    .C(_18413_),
    .Y(_18414_));
 sky130_fd_sc_hd__a21o_2 _28203_ (.A1(_18412_),
    .A2(_18413_),
    .B1(_18411_),
    .X(_18416_));
 sky130_fd_sc_hd__a22o_2 _28204_ (.A1(_17669_),
    .A2(_18164_),
    .B1(_18165_),
    .B2(_18167_),
    .X(_18417_));
 sky130_fd_sc_hd__and3_2 _28205_ (.A(_18414_),
    .B(_18416_),
    .C(_18417_),
    .X(_18418_));
 sky130_fd_sc_hd__a21oi_2 _28206_ (.A1(_18414_),
    .A2(_18416_),
    .B1(_18417_),
    .Y(_18419_));
 sky130_fd_sc_hd__or3_2 _28207_ (.A(_18410_),
    .B(_18418_),
    .C(_18419_),
    .X(_18420_));
 sky130_fd_sc_hd__o21ai_2 _28208_ (.A1(_18418_),
    .A2(_18419_),
    .B1(_18410_),
    .Y(_18421_));
 sky130_fd_sc_hd__and3_2 _28209_ (.A(_18403_),
    .B(_18420_),
    .C(_18421_),
    .X(_18422_));
 sky130_fd_sc_hd__a21oi_2 _28210_ (.A1(_18420_),
    .A2(_18421_),
    .B1(_18403_),
    .Y(_18423_));
 sky130_fd_sc_hd__nor2_2 _28211_ (.A(_18422_),
    .B(_18423_),
    .Y(_18424_));
 sky130_fd_sc_hd__xnor2_2 _28212_ (.A(_18402_),
    .B(_18424_),
    .Y(_18425_));
 sky130_fd_sc_hd__a21oi_2 _28213_ (.A1(_17686_),
    .A2(_18182_),
    .B1(_18184_),
    .Y(_18427_));
 sky130_fd_sc_hd__a31oi_2 _28214_ (.A1(_15887_),
    .A2(_17006_),
    .A3(_18197_),
    .B1(_18195_),
    .Y(_18428_));
 sky130_fd_sc_hd__or3b_2 _28215_ (.A(_12852_),
    .B(_16988_),
    .C_N(_18182_),
    .X(_18429_));
 sky130_fd_sc_hd__a22o_2 _28216_ (.A1(_12846_),
    .A2(_15900_),
    .B1(_16682_),
    .B2(_14634_),
    .X(_18430_));
 sky130_fd_sc_hd__nand2_2 _28217_ (.A(_18429_),
    .B(_18430_),
    .Y(_18431_));
 sky130_fd_sc_hd__nor2_2 _28218_ (.A(_14625_),
    .B(_16312_),
    .Y(_18432_));
 sky130_fd_sc_hd__xor2_2 _28219_ (.A(_18431_),
    .B(_18432_),
    .X(_18433_));
 sky130_fd_sc_hd__xor2_2 _28220_ (.A(_18428_),
    .B(_18433_),
    .X(_18434_));
 sky130_fd_sc_hd__xnor2_2 _28221_ (.A(_18427_),
    .B(_18434_),
    .Y(_18435_));
 sky130_fd_sc_hd__nand2_2 _28222_ (.A(_18192_),
    .B(_17488_),
    .Y(_18436_));
 sky130_fd_sc_hd__and3_2 _28223_ (.A(_12243_),
    .B(_17485_),
    .C(_18194_),
    .X(_18438_));
 sky130_fd_sc_hd__nor2_2 _28224_ (.A(_13926_),
    .B(_17482_),
    .Y(_18439_));
 sky130_fd_sc_hd__a21oi_2 _28225_ (.A1(_14980_),
    .A2(_17702_),
    .B1(_18439_),
    .Y(_18440_));
 sky130_fd_sc_hd__nor2_2 _28226_ (.A(_18438_),
    .B(_18440_),
    .Y(_18441_));
 sky130_fd_sc_hd__xnor2_2 _28227_ (.A(_18436_),
    .B(_18441_),
    .Y(_18442_));
 sky130_fd_sc_hd__nand2_2 _28228_ (.A(_17712_),
    .B(_17713_),
    .Y(_18443_));
 sky130_fd_sc_hd__or3_2 _28229_ (.A(_17708_),
    .B(_17709_),
    .C(_18201_),
    .X(_18444_));
 sky130_fd_sc_hd__or3_2 _28230_ (.A(_16993_),
    .B(_17480_),
    .C(_18444_),
    .X(_18445_));
 sky130_fd_sc_hd__nand2b_2 _28231_ (.A_N(_18445_),
    .B(_16997_),
    .Y(_18446_));
 sky130_fd_sc_hd__nand3b_2 _28232_ (.A_N(_18445_),
    .B(_15663_),
    .C(_16994_),
    .Y(_18447_));
 sky130_fd_sc_hd__a221o_2 _28233_ (.A1(iX[23]),
    .A2(iX[55]),
    .B1(_17706_),
    .B2(_17711_),
    .C1(_17708_),
    .X(_18449_));
 sky130_fd_sc_hd__o21ai_2 _28234_ (.A1(iX[23]),
    .A2(iX[55]),
    .B1(_18449_),
    .Y(_18450_));
 sky130_fd_sc_hd__nand2_2 _28235_ (.A(iX[24]),
    .B(iX[56]),
    .Y(_18451_));
 sky130_fd_sc_hd__or2_2 _28236_ (.A(iX[24]),
    .B(iX[56]),
    .X(_18452_));
 sky130_fd_sc_hd__nand2_2 _28237_ (.A(_18451_),
    .B(_18452_),
    .Y(_18453_));
 sky130_fd_sc_hd__a31o_2 _28238_ (.A1(_18446_),
    .A2(_18447_),
    .A3(_18450_),
    .B1(_18453_),
    .X(_18454_));
 sky130_fd_sc_hd__o211ai_2 _28239_ (.A1(_16998_),
    .A2(_18445_),
    .B1(_18450_),
    .C1(_18453_),
    .Y(_18455_));
 sky130_fd_sc_hd__nand2_2 _28240_ (.A(_18454_),
    .B(_18455_),
    .Y(_18456_));
 sky130_fd_sc_hd__nor2_2 _28241_ (.A(_11576_),
    .B(_18456_),
    .Y(_18457_));
 sky130_fd_sc_hd__and3_2 _28242_ (.A(_11381_),
    .B(_18203_),
    .C(_18457_),
    .X(_18458_));
 sky130_fd_sc_hd__and2_2 _28243_ (.A(_18454_),
    .B(_18455_),
    .X(_18460_));
 sky130_fd_sc_hd__a22o_2 _28244_ (.A1(_11585_),
    .A2(_18203_),
    .B1(_18460_),
    .B2(_11381_),
    .X(_18461_));
 sky130_fd_sc_hd__or4b_4 _28245_ (.A(_11793_),
    .B(_18443_),
    .C(_18458_),
    .D_N(_18461_),
    .X(_18462_));
 sky130_fd_sc_hd__buf_4 _28246_ (.A(_18205_),
    .X(_18463_));
 sky130_fd_sc_hd__or3b_2 _28247_ (.A(_11566_),
    .B(_18210_),
    .C_N(_18457_),
    .X(_18464_));
 sky130_fd_sc_hd__a22o_2 _28248_ (.A1(_15677_),
    .A2(_18463_),
    .B1(_18464_),
    .B2(_18461_),
    .X(_18465_));
 sky130_fd_sc_hd__a31o_2 _28249_ (.A1(_15677_),
    .A2(_18209_),
    .A3(_18206_),
    .B1(_18204_),
    .X(_18466_));
 sky130_fd_sc_hd__nand3_2 _28250_ (.A(_18462_),
    .B(_18465_),
    .C(_18466_),
    .Y(_18467_));
 sky130_fd_sc_hd__a21o_2 _28251_ (.A1(_18462_),
    .A2(_18465_),
    .B1(_18466_),
    .X(_18468_));
 sky130_fd_sc_hd__nand3_2 _28252_ (.A(_18442_),
    .B(_18467_),
    .C(_18468_),
    .Y(_18469_));
 sky130_fd_sc_hd__a21o_4 _28253_ (.A1(_18467_),
    .A2(_18468_),
    .B1(_18442_),
    .X(_18471_));
 sky130_fd_sc_hd__a21bo_4 _28254_ (.A1(_18199_),
    .A2(_18217_),
    .B1_N(_18216_),
    .X(_18472_));
 sky130_fd_sc_hd__nand3_2 _28255_ (.A(_18469_),
    .B(_18471_),
    .C(_18472_),
    .Y(_18473_));
 sky130_fd_sc_hd__a21o_4 _28256_ (.A1(_18469_),
    .A2(_18471_),
    .B1(_18472_),
    .X(_18474_));
 sky130_fd_sc_hd__nand3_2 _28257_ (.A(_18435_),
    .B(_18473_),
    .C(_18474_),
    .Y(_18475_));
 sky130_fd_sc_hd__a21o_4 _28258_ (.A1(_18473_),
    .A2(_18474_),
    .B1(_18435_),
    .X(_18476_));
 sky130_fd_sc_hd__o211ai_2 _28259_ (.A1(_18223_),
    .A2(_18225_),
    .B1(_18475_),
    .C1(_18476_),
    .Y(_18477_));
 sky130_fd_sc_hd__a211o_2 _28260_ (.A1(_18475_),
    .A2(_18476_),
    .B1(_18223_),
    .C1(_18225_),
    .X(_18478_));
 sky130_fd_sc_hd__and3_4 _28261_ (.A(_18425_),
    .B(_18477_),
    .C(_18478_),
    .X(_18479_));
 sky130_fd_sc_hd__a21oi_2 _28262_ (.A1(_18477_),
    .A2(_18478_),
    .B1(_18425_),
    .Y(_18480_));
 sky130_fd_sc_hd__a211o_4 _28263_ (.A1(_18227_),
    .A2(_18401_),
    .B1(_18479_),
    .C1(_18480_),
    .X(_18482_));
 sky130_fd_sc_hd__o211ai_2 _28264_ (.A1(_18479_),
    .A2(_18480_),
    .B1(_18227_),
    .C1(_18401_),
    .Y(_18483_));
 sky130_fd_sc_hd__nand3_2 _28265_ (.A(_18400_),
    .B(_18482_),
    .C(_18483_),
    .Y(_18484_));
 sky130_fd_sc_hd__a21o_2 _28266_ (.A1(_18482_),
    .A2(_18483_),
    .B1(_18400_),
    .X(_18485_));
 sky130_fd_sc_hd__o211ai_2 _28267_ (.A1(_18232_),
    .A2(_18234_),
    .B1(_18484_),
    .C1(_18485_),
    .Y(_18486_));
 sky130_fd_sc_hd__a211o_4 _28268_ (.A1(_18484_),
    .A2(_18485_),
    .B1(_18232_),
    .C1(_18234_),
    .X(_18487_));
 sky130_fd_sc_hd__nand3_2 _28269_ (.A(_18354_),
    .B(_18486_),
    .C(_18487_),
    .Y(_18488_));
 sky130_fd_sc_hd__a21o_4 _28270_ (.A1(_18486_),
    .A2(_18487_),
    .B1(_18354_),
    .X(_18489_));
 sky130_fd_sc_hd__o211ai_2 _28271_ (.A1(_18323_),
    .A2(_18238_),
    .B1(_18488_),
    .C1(_18489_),
    .Y(_18490_));
 sky130_fd_sc_hd__a211o_2 _28272_ (.A1(_18488_),
    .A2(_18489_),
    .B1(_18323_),
    .C1(_18238_),
    .X(_18491_));
 sky130_fd_sc_hd__nand3_2 _28273_ (.A(_18322_),
    .B(_18490_),
    .C(_18491_),
    .Y(_18493_));
 sky130_fd_sc_hd__a21o_2 _28274_ (.A1(_18490_),
    .A2(_18491_),
    .B1(_18322_),
    .X(_18494_));
 sky130_fd_sc_hd__o211a_2 _28275_ (.A1(_18320_),
    .A2(_18321_),
    .B1(_18493_),
    .C1(_18494_),
    .X(_18495_));
 sky130_fd_sc_hd__a211oi_2 _28276_ (.A1(_18493_),
    .A2(_18494_),
    .B1(_18320_),
    .C1(_18321_),
    .Y(_18496_));
 sky130_fd_sc_hd__nor3_2 _28277_ (.A(_18245_),
    .B(_18495_),
    .C(_18496_),
    .Y(_18497_));
 sky130_fd_sc_hd__o21a_2 _28278_ (.A1(_18495_),
    .A2(_18496_),
    .B1(_18245_),
    .X(_18498_));
 sky130_fd_sc_hd__or2_2 _28279_ (.A(_18497_),
    .B(_18498_),
    .X(_18499_));
 sky130_fd_sc_hd__xnor2_2 _28280_ (.A(_18319_),
    .B(_18499_),
    .Y(_18500_));
 sky130_fd_sc_hd__a21oi_2 _28281_ (.A1(_17260_),
    .A2(_17372_),
    .B1(_17866_),
    .Y(_18501_));
 sky130_fd_sc_hd__or3_2 _28282_ (.A(_17865_),
    .B(_18501_),
    .C(_18077_),
    .X(_18502_));
 sky130_fd_sc_hd__a21o_2 _28283_ (.A1(_17948_),
    .A2(_18078_),
    .B1(_18076_),
    .X(_18504_));
 sky130_fd_sc_hd__inv_2 _28284_ (.A(_17372_),
    .Y(_18505_));
 sky130_fd_sc_hd__or4_2 _28285_ (.A(_17162_),
    .B(_18505_),
    .C(_17865_),
    .D(_18077_),
    .X(_18506_));
 sky130_fd_sc_hd__a211o_2 _28286_ (.A1(_17163_),
    .A2(_17165_),
    .B1(_17167_),
    .C1(_18506_),
    .X(_18507_));
 sky130_fd_sc_hd__nand3_2 _28287_ (.A(_18502_),
    .B(_18504_),
    .C(_18507_),
    .Y(_18508_));
 sky130_fd_sc_hd__or2_2 _28288_ (.A(_18072_),
    .B(_18074_),
    .X(_18509_));
 sky130_fd_sc_hd__nand2_2 _28289_ (.A(_18059_),
    .B(_18065_),
    .Y(_18510_));
 sky130_fd_sc_hd__nand3_2 _28290_ (.A(_18011_),
    .B(_18012_),
    .C(_18052_),
    .Y(_18511_));
 sky130_fd_sc_hd__and3_2 _28291_ (.A(_17979_),
    .B(_17980_),
    .C(_17982_),
    .X(_18512_));
 sky130_fd_sc_hd__or2b_2 _28292_ (.A(_17958_),
    .B_N(_17957_),
    .X(_18513_));
 sky130_fd_sc_hd__nand2_2 _28293_ (.A(_17959_),
    .B(_17964_),
    .Y(_18515_));
 sky130_fd_sc_hd__and4_2 _28294_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[53]),
    .D(iX[54]),
    .X(_18516_));
 sky130_fd_sc_hd__a22oi_2 _28295_ (.A1(iY[35]),
    .A2(iX[53]),
    .B1(iX[54]),
    .B2(iY[34]),
    .Y(_18517_));
 sky130_fd_sc_hd__nor2_2 _28296_ (.A(_18516_),
    .B(_18517_),
    .Y(_18518_));
 sky130_fd_sc_hd__nand2_2 _28297_ (.A(iY[33]),
    .B(iX[55]),
    .Y(_18519_));
 sky130_fd_sc_hd__xnor2_2 _28298_ (.A(_18518_),
    .B(_18519_),
    .Y(_18520_));
 sky130_fd_sc_hd__o21ba_2 _28299_ (.A1(_17953_),
    .A2(_17956_),
    .B1_N(_17952_),
    .X(_18521_));
 sky130_fd_sc_hd__xnor2_2 _28300_ (.A(_18520_),
    .B(_18521_),
    .Y(_18522_));
 sky130_fd_sc_hd__and4_2 _28301_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[52]),
    .D(iX[56]),
    .X(_18523_));
 sky130_fd_sc_hd__a22oi_2 _28302_ (.A1(iY[36]),
    .A2(iX[52]),
    .B1(iX[56]),
    .B2(iY[32]),
    .Y(_18524_));
 sky130_fd_sc_hd__nor2_2 _28303_ (.A(_18523_),
    .B(_18524_),
    .Y(_18526_));
 sky130_fd_sc_hd__nand2_2 _28304_ (.A(iY[37]),
    .B(iX[51]),
    .Y(_18527_));
 sky130_fd_sc_hd__xnor2_2 _28305_ (.A(_18526_),
    .B(_18527_),
    .Y(_18528_));
 sky130_fd_sc_hd__xnor2_2 _28306_ (.A(_18522_),
    .B(_18528_),
    .Y(_18529_));
 sky130_fd_sc_hd__a21o_2 _28307_ (.A1(_18513_),
    .A2(_18515_),
    .B1(_18529_),
    .X(_18530_));
 sky130_fd_sc_hd__nand3_2 _28308_ (.A(_18513_),
    .B(_18515_),
    .C(_18529_),
    .Y(_18531_));
 sky130_fd_sc_hd__o21ba_2 _28309_ (.A1(_17972_),
    .A2(_17974_),
    .B1_N(_17971_),
    .X(_18532_));
 sky130_fd_sc_hd__o21ba_2 _28310_ (.A1(_17961_),
    .A2(_17963_),
    .B1_N(_17960_),
    .X(_18533_));
 sky130_fd_sc_hd__and4_2 _28311_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[49]),
    .D(iX[50]),
    .X(_18534_));
 sky130_fd_sc_hd__a22oi_2 _28312_ (.A1(iY[39]),
    .A2(iX[49]),
    .B1(iX[50]),
    .B2(iY[38]),
    .Y(_18535_));
 sky130_fd_sc_hd__nor2_2 _28313_ (.A(_18534_),
    .B(_18535_),
    .Y(_18537_));
 sky130_fd_sc_hd__nand2_2 _28314_ (.A(iY[40]),
    .B(iX[48]),
    .Y(_18538_));
 sky130_fd_sc_hd__xnor2_2 _28315_ (.A(_18537_),
    .B(_18538_),
    .Y(_18539_));
 sky130_fd_sc_hd__xnor2_2 _28316_ (.A(_18533_),
    .B(_18539_),
    .Y(_18540_));
 sky130_fd_sc_hd__xnor2_2 _28317_ (.A(_18532_),
    .B(_18540_),
    .Y(_18541_));
 sky130_fd_sc_hd__and3_2 _28318_ (.A(_18530_),
    .B(_18531_),
    .C(_18541_),
    .X(_18542_));
 sky130_fd_sc_hd__a21oi_2 _28319_ (.A1(_18530_),
    .A2(_18531_),
    .B1(_18541_),
    .Y(_18543_));
 sky130_fd_sc_hd__nor2_2 _28320_ (.A(_18542_),
    .B(_18543_),
    .Y(_18544_));
 sky130_fd_sc_hd__nand2_2 _28321_ (.A(_17967_),
    .B(_17979_),
    .Y(_18545_));
 sky130_fd_sc_hd__xnor2_2 _28322_ (.A(_18544_),
    .B(_18545_),
    .Y(_18546_));
 sky130_fd_sc_hd__and2b_2 _28323_ (.A_N(_17999_),
    .B(_17997_),
    .X(_18548_));
 sky130_fd_sc_hd__or2b_2 _28324_ (.A(_17970_),
    .B_N(_17975_),
    .X(_18549_));
 sky130_fd_sc_hd__or2b_2 _28325_ (.A(_17969_),
    .B_N(_17977_),
    .X(_18550_));
 sky130_fd_sc_hd__and4_2 _28326_ (.A(iX[43]),
    .B(iX[44]),
    .C(iY[44]),
    .D(iY[45]),
    .X(_18551_));
 sky130_fd_sc_hd__a22oi_2 _28327_ (.A1(iX[44]),
    .A2(iY[44]),
    .B1(iY[45]),
    .B2(iX[43]),
    .Y(_18552_));
 sky130_fd_sc_hd__nor2_2 _28328_ (.A(_18551_),
    .B(_18552_),
    .Y(_18553_));
 sky130_fd_sc_hd__nand2_2 _28329_ (.A(iX[42]),
    .B(iY[46]),
    .Y(_18554_));
 sky130_fd_sc_hd__xnor2_2 _28330_ (.A(_18553_),
    .B(_18554_),
    .Y(_18555_));
 sky130_fd_sc_hd__and4_2 _28331_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[46]),
    .D(iX[47]),
    .X(_18556_));
 sky130_fd_sc_hd__a22oi_2 _28332_ (.A1(iY[42]),
    .A2(iX[46]),
    .B1(iX[47]),
    .B2(iY[41]),
    .Y(_18557_));
 sky130_fd_sc_hd__nor2_2 _28333_ (.A(_18556_),
    .B(_18557_),
    .Y(_18559_));
 sky130_fd_sc_hd__nand2_2 _28334_ (.A(iY[43]),
    .B(iX[45]),
    .Y(_18560_));
 sky130_fd_sc_hd__xnor2_2 _28335_ (.A(_18559_),
    .B(_18560_),
    .Y(_18561_));
 sky130_fd_sc_hd__nor2_2 _28336_ (.A(_17993_),
    .B(_17995_),
    .Y(_18562_));
 sky130_fd_sc_hd__xnor2_2 _28337_ (.A(_18561_),
    .B(_18562_),
    .Y(_18563_));
 sky130_fd_sc_hd__xnor2_2 _28338_ (.A(_18555_),
    .B(_18563_),
    .Y(_18564_));
 sky130_fd_sc_hd__a21oi_2 _28339_ (.A1(_18549_),
    .A2(_18550_),
    .B1(_18564_),
    .Y(_18565_));
 sky130_fd_sc_hd__inv_2 _28340_ (.A(_18565_),
    .Y(_18566_));
 sky130_fd_sc_hd__nand3_2 _28341_ (.A(_18549_),
    .B(_18550_),
    .C(_18564_),
    .Y(_18567_));
 sky130_fd_sc_hd__o211a_2 _28342_ (.A1(_18548_),
    .A2(_18001_),
    .B1(_18566_),
    .C1(_18567_),
    .X(_18568_));
 sky130_fd_sc_hd__a211o_2 _28343_ (.A1(_18566_),
    .A2(_18567_),
    .B1(_18548_),
    .C1(_18001_),
    .X(_18570_));
 sky130_fd_sc_hd__or3b_2 _28344_ (.A(_18546_),
    .B(_18568_),
    .C_N(_18570_),
    .X(_18571_));
 sky130_fd_sc_hd__inv_2 _28345_ (.A(_18568_),
    .Y(_18572_));
 sky130_fd_sc_hd__a21bo_2 _28346_ (.A1(_18572_),
    .A2(_18570_),
    .B1_N(_18546_),
    .X(_18573_));
 sky130_fd_sc_hd__o211a_2 _28347_ (.A1(_18512_),
    .A2(_18008_),
    .B1(_18571_),
    .C1(_18573_),
    .X(_18574_));
 sky130_fd_sc_hd__a211oi_2 _28348_ (.A1(_18571_),
    .A2(_18573_),
    .B1(_18512_),
    .C1(_18008_),
    .Y(_18575_));
 sky130_fd_sc_hd__inv_2 _28349_ (.A(_18043_),
    .Y(_18576_));
 sky130_fd_sc_hd__and4_2 _28350_ (.A(iX[34]),
    .B(iX[35]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_18577_));
 sky130_fd_sc_hd__a22oi_2 _28351_ (.A1(iX[35]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[34]),
    .Y(_18578_));
 sky130_fd_sc_hd__nor2_2 _28352_ (.A(_18577_),
    .B(_18578_),
    .Y(_18579_));
 sky130_fd_sc_hd__nand2_2 _28353_ (.A(iX[33]),
    .B(iY[55]),
    .Y(_18581_));
 sky130_fd_sc_hd__xnor2_2 _28354_ (.A(_18579_),
    .B(_18581_),
    .Y(_18582_));
 sky130_fd_sc_hd__and4_2 _28355_ (.A(iX[37]),
    .B(iX[38]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_18583_));
 sky130_fd_sc_hd__a22oi_2 _28356_ (.A1(iX[38]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[37]),
    .Y(_18584_));
 sky130_fd_sc_hd__nor2_2 _28357_ (.A(_18583_),
    .B(_18584_),
    .Y(_18585_));
 sky130_fd_sc_hd__nand2_2 _28358_ (.A(iX[36]),
    .B(iY[52]),
    .Y(_18586_));
 sky130_fd_sc_hd__xnor2_2 _28359_ (.A(_18585_),
    .B(_18586_),
    .Y(_18587_));
 sky130_fd_sc_hd__a31o_2 _28360_ (.A1(iX[35]),
    .A2(iY[52]),
    .A3(_18021_),
    .B1(_18019_),
    .X(_18588_));
 sky130_fd_sc_hd__xor2_2 _28361_ (.A(_18587_),
    .B(_18588_),
    .X(_18589_));
 sky130_fd_sc_hd__and2_2 _28362_ (.A(_18582_),
    .B(_18589_),
    .X(_18590_));
 sky130_fd_sc_hd__nor2_2 _28363_ (.A(_18582_),
    .B(_18589_),
    .Y(_18592_));
 sky130_fd_sc_hd__or2_2 _28364_ (.A(_18590_),
    .B(_18592_),
    .X(_18593_));
 sky130_fd_sc_hd__or3_2 _28365_ (.A(_18034_),
    .B(_18037_),
    .C(_18038_),
    .X(_18594_));
 sky130_fd_sc_hd__nand2_2 _28366_ (.A(_18033_),
    .B(_18040_),
    .Y(_18595_));
 sky130_fd_sc_hd__o21ba_2 _28367_ (.A1(_17989_),
    .A2(_17991_),
    .B1_N(_17988_),
    .X(_18596_));
 sky130_fd_sc_hd__and4_2 _28368_ (.A(iX[40]),
    .B(iX[41]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_18597_));
 sky130_fd_sc_hd__a22oi_2 _28369_ (.A1(iX[41]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[40]),
    .Y(_18598_));
 sky130_fd_sc_hd__and4bb_2 _28370_ (.A_N(_18597_),
    .B_N(_18598_),
    .C(iX[39]),
    .D(iY[49]),
    .X(_18599_));
 sky130_fd_sc_hd__o2bb2a_2 _28371_ (.A1_N(iX[39]),
    .A2_N(iY[49]),
    .B1(_18597_),
    .B2(_18598_),
    .X(_18600_));
 sky130_fd_sc_hd__nor2_2 _28372_ (.A(_18599_),
    .B(_18600_),
    .Y(_18601_));
 sky130_fd_sc_hd__xnor2_2 _28373_ (.A(_18596_),
    .B(_18601_),
    .Y(_18603_));
 sky130_fd_sc_hd__o21ai_2 _28374_ (.A1(_18035_),
    .A2(_18037_),
    .B1(_18603_),
    .Y(_18604_));
 sky130_fd_sc_hd__or3_2 _28375_ (.A(_18035_),
    .B(_18037_),
    .C(_18603_),
    .X(_18605_));
 sky130_fd_sc_hd__nand2_2 _28376_ (.A(_18604_),
    .B(_18605_),
    .Y(_18606_));
 sky130_fd_sc_hd__a21oi_2 _28377_ (.A1(_18594_),
    .A2(_18595_),
    .B1(_18606_),
    .Y(_18607_));
 sky130_fd_sc_hd__and3_2 _28378_ (.A(_18594_),
    .B(_18595_),
    .C(_18606_),
    .X(_18608_));
 sky130_fd_sc_hd__nor3_2 _28379_ (.A(_18593_),
    .B(_18607_),
    .C(_18608_),
    .Y(_18609_));
 sky130_fd_sc_hd__o21a_2 _28380_ (.A1(_18607_),
    .A2(_18608_),
    .B1(_18593_),
    .X(_18610_));
 sky130_fd_sc_hd__a211oi_2 _28381_ (.A1(_18004_),
    .A2(_18006_),
    .B1(_18609_),
    .C1(_18610_),
    .Y(_18611_));
 sky130_fd_sc_hd__o211a_2 _28382_ (.A1(_18609_),
    .A2(_18610_),
    .B1(_18004_),
    .C1(_18006_),
    .X(_18612_));
 sky130_fd_sc_hd__a211oi_2 _28383_ (.A1(_18576_),
    .A2(_18045_),
    .B1(_18611_),
    .C1(_18612_),
    .Y(_18614_));
 sky130_fd_sc_hd__o211a_2 _28384_ (.A1(_18611_),
    .A2(_18612_),
    .B1(_18576_),
    .C1(_18045_),
    .X(_18615_));
 sky130_fd_sc_hd__nor4_2 _28385_ (.A(_18574_),
    .B(_18575_),
    .C(_18614_),
    .D(_18615_),
    .Y(_18616_));
 sky130_fd_sc_hd__o22a_2 _28386_ (.A1(_18574_),
    .A2(_18575_),
    .B1(_18614_),
    .B2(_18615_),
    .X(_18617_));
 sky130_fd_sc_hd__a211oi_2 _28387_ (.A1(_18011_),
    .A2(_18511_),
    .B1(_18616_),
    .C1(_18617_),
    .Y(_18618_));
 sky130_fd_sc_hd__o211a_2 _28388_ (.A1(_18616_),
    .A2(_18617_),
    .B1(_18011_),
    .C1(_18511_),
    .X(_18619_));
 sky130_fd_sc_hd__or2_2 _28389_ (.A(_18618_),
    .B(_18619_),
    .X(_18620_));
 sky130_fd_sc_hd__and2_2 _28390_ (.A(_18024_),
    .B(_18025_),
    .X(_18621_));
 sky130_fd_sc_hd__a31o_2 _28391_ (.A1(iX[32]),
    .A2(iY[55]),
    .A3(_18015_),
    .B1(_18014_),
    .X(_18622_));
 sky130_fd_sc_hd__and3_2 _28392_ (.A(iX[32]),
    .B(iY[56]),
    .C(_18622_),
    .X(_18623_));
 sky130_fd_sc_hd__a21oi_2 _28393_ (.A1(iX[32]),
    .A2(iY[56]),
    .B1(_18622_),
    .Y(_18625_));
 sky130_fd_sc_hd__nor2_2 _28394_ (.A(_18623_),
    .B(_18625_),
    .Y(_18626_));
 sky130_fd_sc_hd__o21ai_2 _28395_ (.A1(_18621_),
    .A2(_18027_),
    .B1(_18626_),
    .Y(_18627_));
 sky130_fd_sc_hd__or3_2 _28396_ (.A(_18621_),
    .B(_18027_),
    .C(_18626_),
    .X(_18628_));
 sky130_fd_sc_hd__and2_2 _28397_ (.A(_18627_),
    .B(_18628_),
    .X(_18629_));
 sky130_fd_sc_hd__xnor2_2 _28398_ (.A(_18062_),
    .B(_18629_),
    .Y(_18630_));
 sky130_fd_sc_hd__o21a_2 _28399_ (.A1(_18048_),
    .A2(_18050_),
    .B1(_18630_),
    .X(_18631_));
 sky130_fd_sc_hd__nor3_2 _28400_ (.A(_18048_),
    .B(_18050_),
    .C(_18630_),
    .Y(_18632_));
 sky130_fd_sc_hd__or2_2 _28401_ (.A(_18631_),
    .B(_18632_),
    .X(_18633_));
 sky130_fd_sc_hd__nor2_2 _28402_ (.A(_18620_),
    .B(_18633_),
    .Y(_18634_));
 sky130_fd_sc_hd__and2_2 _28403_ (.A(_18620_),
    .B(_18633_),
    .X(_18636_));
 sky130_fd_sc_hd__or2_2 _28404_ (.A(_18634_),
    .B(_18636_),
    .X(_18637_));
 sky130_fd_sc_hd__o31a_2 _28405_ (.A1(_18054_),
    .A2(_18055_),
    .A3(_18057_),
    .B1(_18067_),
    .X(_18638_));
 sky130_fd_sc_hd__xnor2_2 _28406_ (.A(_18637_),
    .B(_18638_),
    .Y(_18639_));
 sky130_fd_sc_hd__xor2_2 _28407_ (.A(_18510_),
    .B(_18639_),
    .X(_18640_));
 sky130_fd_sc_hd__a32o_2 _28408_ (.A1(_18067_),
    .A2(_18068_),
    .A3(_18070_),
    .B1(_18071_),
    .B2(_17854_),
    .X(_18641_));
 sky130_fd_sc_hd__xnor2_2 _28409_ (.A(_18640_),
    .B(_18641_),
    .Y(_18642_));
 sky130_fd_sc_hd__nor2_2 _28410_ (.A(_18509_),
    .B(_18642_),
    .Y(_18643_));
 sky130_fd_sc_hd__and2_2 _28411_ (.A(_18509_),
    .B(_18642_),
    .X(_18644_));
 sky130_fd_sc_hd__nor2_2 _28412_ (.A(_18643_),
    .B(_18644_),
    .Y(_18645_));
 sky130_fd_sc_hd__xor2_2 _28413_ (.A(_18508_),
    .B(_18645_),
    .X(_18647_));
 sky130_fd_sc_hd__xnor2_2 _28414_ (.A(_18500_),
    .B(_18647_),
    .Y(_18648_));
 sky130_fd_sc_hd__xnor2_2 _28415_ (.A(_09530_),
    .B(_18648_),
    .Y(_18649_));
 sky130_fd_sc_hd__and2b_2 _28416_ (.A_N(_18256_),
    .B(_18080_),
    .X(_18650_));
 sky130_fd_sc_hd__a21oi_2 _28417_ (.A1(_08066_),
    .A2(_18257_),
    .B1(_18650_),
    .Y(_18651_));
 sky130_fd_sc_hd__xnor2_2 _28418_ (.A(_18649_),
    .B(_18651_),
    .Y(_18652_));
 sky130_fd_sc_hd__a21o_2 _28419_ (.A1(_17946_),
    .A2(_17947_),
    .B1(_18258_),
    .X(_18653_));
 sky130_fd_sc_hd__o211a_2 _28420_ (.A1(_17873_),
    .A2(_18259_),
    .B1(_18653_),
    .C1(_17880_),
    .X(_18654_));
 sky130_fd_sc_hd__nor2_2 _28421_ (.A(_17874_),
    .B(_18260_),
    .Y(_18655_));
 sky130_fd_sc_hd__a211o_2 _28422_ (.A1(_17877_),
    .A2(_18654_),
    .B1(_18655_),
    .C1(_18259_),
    .X(_18656_));
 sky130_fd_sc_hd__xor2_2 _28423_ (.A(_18652_),
    .B(_18656_),
    .X(_18658_));
 sky130_fd_sc_hd__xor2_2 _28424_ (.A(_18312_),
    .B(_18658_),
    .X(_18659_));
 sky130_fd_sc_hd__inv_2 _28425_ (.A(_18659_),
    .Y(_18660_));
 sky130_fd_sc_hd__nand2_2 _28426_ (.A(_17944_),
    .B(_18263_),
    .Y(_18661_));
 sky130_fd_sc_hd__nor2_2 _28427_ (.A(_17944_),
    .B(_18263_),
    .Y(_18662_));
 sky130_fd_sc_hd__nand2_2 _28428_ (.A(_17885_),
    .B(_18264_),
    .Y(_18663_));
 sky130_fd_sc_hd__nor2_2 _28429_ (.A(_17887_),
    .B(_18663_),
    .Y(_18664_));
 sky130_fd_sc_hd__a211o_2 _28430_ (.A1(_17883_),
    .A2(_18661_),
    .B1(_18662_),
    .C1(_18664_),
    .X(_18665_));
 sky130_fd_sc_hd__or4b_2 _28431_ (.A(_17184_),
    .B(_18663_),
    .C(_17535_),
    .D_N(_17886_),
    .X(_18666_));
 sky130_fd_sc_hd__a221oi_2 _28432_ (.A1(_16481_),
    .A2(_17187_),
    .B1(_17189_),
    .B2(_17186_),
    .C1(_18666_),
    .Y(_18667_));
 sky130_fd_sc_hd__nor2_2 _28433_ (.A(_18665_),
    .B(_18667_),
    .Y(_18669_));
 sky130_fd_sc_hd__xnor2_2 _28434_ (.A(_18660_),
    .B(_18669_),
    .Y(oO[56]));
 sky130_fd_sc_hd__nand2_2 _28435_ (.A(_18270_),
    .B(_18311_),
    .Y(_18670_));
 sky130_fd_sc_hd__or2b_2 _28436_ (.A(_18279_),
    .B_N(_18278_),
    .X(_18671_));
 sky130_fd_sc_hd__and4_2 _28437_ (.A(iY[27]),
    .B(iY[28]),
    .C(iX[29]),
    .D(iX[30]),
    .X(_18672_));
 sky130_fd_sc_hd__a22oi_2 _28438_ (.A1(iY[28]),
    .A2(iX[29]),
    .B1(iX[30]),
    .B2(iY[27]),
    .Y(_18673_));
 sky130_fd_sc_hd__nor2_2 _28439_ (.A(_18672_),
    .B(_18673_),
    .Y(_18674_));
 sky130_fd_sc_hd__nand2_2 _28440_ (.A(iX[28]),
    .B(iY[29]),
    .Y(_18675_));
 sky130_fd_sc_hd__xnor2_2 _28441_ (.A(_18674_),
    .B(_18675_),
    .Y(_18676_));
 sky130_fd_sc_hd__o21ba_2 _28442_ (.A1(_18275_),
    .A2(_18277_),
    .B1_N(_18274_),
    .X(_18677_));
 sky130_fd_sc_hd__xnor2_2 _28443_ (.A(_18676_),
    .B(_18677_),
    .Y(_18679_));
 sky130_fd_sc_hd__nand3_2 _28444_ (.A(iX[27]),
    .B(iY[30]),
    .C(_18679_),
    .Y(_18680_));
 sky130_fd_sc_hd__a21o_2 _28445_ (.A1(iX[27]),
    .A2(iY[30]),
    .B1(_18679_),
    .X(_18681_));
 sky130_fd_sc_hd__nand2_2 _28446_ (.A(_18680_),
    .B(_18681_),
    .Y(_18682_));
 sky130_fd_sc_hd__a21o_2 _28447_ (.A1(_18671_),
    .A2(_18281_),
    .B1(_18682_),
    .X(_18683_));
 sky130_fd_sc_hd__nand3_2 _28448_ (.A(_18671_),
    .B(_18281_),
    .C(_18682_),
    .Y(_18684_));
 sky130_fd_sc_hd__and2_2 _28449_ (.A(_18683_),
    .B(_18684_),
    .X(_18685_));
 sky130_fd_sc_hd__a21o_2 _28450_ (.A1(iX[26]),
    .A2(iY[31]),
    .B1(_18685_),
    .X(_18686_));
 sky130_fd_sc_hd__nand3_2 _28451_ (.A(iX[26]),
    .B(iY[31]),
    .C(_18685_),
    .Y(_18687_));
 sky130_fd_sc_hd__and2_2 _28452_ (.A(_18686_),
    .B(_18687_),
    .X(_18688_));
 sky130_fd_sc_hd__and3b_2 _28453_ (.A_N(_17543_),
    .B(iX[31]),
    .C(iY[26]),
    .X(_18690_));
 sky130_fd_sc_hd__and3_2 _28454_ (.A(_17896_),
    .B(_17897_),
    .C(_18298_),
    .X(_18691_));
 sky130_fd_sc_hd__nor2_2 _28455_ (.A(_18296_),
    .B(_18691_),
    .Y(_18692_));
 sky130_fd_sc_hd__xnor2_2 _28456_ (.A(_18690_),
    .B(_18692_),
    .Y(_18693_));
 sky130_fd_sc_hd__xor2_2 _28457_ (.A(_18688_),
    .B(_18693_),
    .X(_18694_));
 sky130_fd_sc_hd__a22o_2 _28458_ (.A1(_17901_),
    .A2(_18298_),
    .B1(_18300_),
    .B2(_18290_),
    .X(_18695_));
 sky130_fd_sc_hd__and2_2 _28459_ (.A(_18694_),
    .B(_18695_),
    .X(_18696_));
 sky130_fd_sc_hd__nor2_2 _28460_ (.A(_18694_),
    .B(_18695_),
    .Y(_18697_));
 sky130_fd_sc_hd__nor2_2 _28461_ (.A(_18696_),
    .B(_18697_),
    .Y(_18698_));
 sky130_fd_sc_hd__and3b_2 _28462_ (.A_N(_18302_),
    .B(_18303_),
    .C(_17928_),
    .X(_18699_));
 sky130_fd_sc_hd__or2_2 _28463_ (.A(_18302_),
    .B(_18699_),
    .X(_18701_));
 sky130_fd_sc_hd__xnor2_2 _28464_ (.A(_18698_),
    .B(_18701_),
    .Y(_18702_));
 sky130_fd_sc_hd__a21oi_2 _28465_ (.A1(_18285_),
    .A2(_18289_),
    .B1(_18702_),
    .Y(_18703_));
 sky130_fd_sc_hd__and3_2 _28466_ (.A(_18285_),
    .B(_18289_),
    .C(_18702_),
    .X(_18704_));
 sky130_fd_sc_hd__nor2_2 _28467_ (.A(_18703_),
    .B(_18704_),
    .Y(_18705_));
 sky130_fd_sc_hd__inv_2 _28468_ (.A(_18705_),
    .Y(_18706_));
 sky130_fd_sc_hd__a32oi_2 _28469_ (.A1(_17930_),
    .A2(_17931_),
    .A3(_18306_),
    .B1(_18307_),
    .B2(_18308_),
    .Y(_18707_));
 sky130_fd_sc_hd__xnor2_2 _28470_ (.A(_18706_),
    .B(_18707_),
    .Y(_18708_));
 sky130_fd_sc_hd__inv_2 _28471_ (.A(_18708_),
    .Y(_18709_));
 sky130_fd_sc_hd__and2b_2 _28472_ (.A_N(_18309_),
    .B(_18310_),
    .X(_18710_));
 sky130_fd_sc_hd__a211o_2 _28473_ (.A1(_18270_),
    .A2(_18311_),
    .B1(_18709_),
    .C1(_18710_),
    .X(_18712_));
 sky130_fd_sc_hd__nand2_2 _28474_ (.A(_18710_),
    .B(_18709_),
    .Y(_18713_));
 sky130_fd_sc_hd__o211ai_2 _28475_ (.A1(_18670_),
    .A2(_18708_),
    .B1(_18712_),
    .C1(_18713_),
    .Y(_18714_));
 sky130_fd_sc_hd__or3_2 _28476_ (.A(_18245_),
    .B(_18495_),
    .C(_18496_),
    .X(_18715_));
 sky130_fd_sc_hd__a21o_2 _28477_ (.A1(_18315_),
    .A2(_18318_),
    .B1(_18499_),
    .X(_18716_));
 sky130_fd_sc_hd__a21oi_2 _28478_ (.A1(_18355_),
    .A2(_18399_),
    .B1(_18397_),
    .Y(_18717_));
 sky130_fd_sc_hd__or2b_2 _28479_ (.A(_18346_),
    .B_N(_18325_),
    .X(_18718_));
 sky130_fd_sc_hd__and2_2 _28480_ (.A(_18330_),
    .B(_18345_),
    .X(_18719_));
 sky130_fd_sc_hd__nand2_2 _28481_ (.A(_18374_),
    .B(_18376_),
    .Y(_18720_));
 sky130_fd_sc_hd__nor2_2 _28482_ (.A(_18100_),
    .B(_18358_),
    .Y(_18721_));
 sky130_fd_sc_hd__a31o_2 _28483_ (.A1(_17392_),
    .A2(_18326_),
    .A3(_18359_),
    .B1(_18721_),
    .X(_18723_));
 sky130_fd_sc_hd__nor2_2 _28484_ (.A(iY[25]),
    .B(iY[57]),
    .Y(_18724_));
 sky130_fd_sc_hd__and2_2 _28485_ (.A(iY[25]),
    .B(iY[57]),
    .X(_18725_));
 sky130_fd_sc_hd__or2_2 _28486_ (.A(_18724_),
    .B(_18725_),
    .X(_18726_));
 sky130_fd_sc_hd__o31a_2 _28487_ (.A1(_18333_),
    .A2(_18337_),
    .A3(_18339_),
    .B1(_18331_),
    .X(_18727_));
 sky130_fd_sc_hd__xor2_2 _28488_ (.A(_18726_),
    .B(_18727_),
    .X(_18728_));
 sky130_fd_sc_hd__buf_2 _28489_ (.A(_18728_),
    .X(_18729_));
 sky130_fd_sc_hd__o2bb2a_2 _28490_ (.A1_N(_14592_),
    .A2_N(_18729_),
    .B1(_18343_),
    .B2(_11571_),
    .X(_18730_));
 sky130_fd_sc_hd__and2_4 _28491_ (.A(_18340_),
    .B(_18341_),
    .X(_18731_));
 sky130_fd_sc_hd__buf_2 _28492_ (.A(_18731_),
    .X(_18732_));
 sky130_fd_sc_hd__buf_4 _28493_ (.A(_18732_),
    .X(_18734_));
 sky130_fd_sc_hd__and4_2 _28494_ (.A(_14592_),
    .B(_17392_),
    .C(_18734_),
    .D(_18729_),
    .X(_18735_));
 sky130_fd_sc_hd__nor2_2 _28495_ (.A(_18730_),
    .B(_18735_),
    .Y(_18736_));
 sky130_fd_sc_hd__nand2_2 _28496_ (.A(_18723_),
    .B(_18736_),
    .Y(_18737_));
 sky130_fd_sc_hd__or2_2 _28497_ (.A(_18723_),
    .B(_18736_),
    .X(_18738_));
 sky130_fd_sc_hd__nand2_2 _28498_ (.A(_18737_),
    .B(_18738_),
    .Y(_18739_));
 sky130_fd_sc_hd__xnor2_2 _28499_ (.A(_18720_),
    .B(_18739_),
    .Y(_18740_));
 sky130_fd_sc_hd__xnor2_2 _28500_ (.A(_18719_),
    .B(_18740_),
    .Y(_18741_));
 sky130_fd_sc_hd__xor2_2 _28501_ (.A(_18718_),
    .B(_18741_),
    .X(_18742_));
 sky130_fd_sc_hd__xnor2_2 _28502_ (.A(_18717_),
    .B(_18742_),
    .Y(_18743_));
 sky130_fd_sc_hd__xnor2_2 _28503_ (.A(_18348_),
    .B(_18743_),
    .Y(_18745_));
 sky130_fd_sc_hd__nand2_2 _28504_ (.A(_18392_),
    .B(_18395_),
    .Y(_18746_));
 sky130_fd_sc_hd__o21bai_2 _28505_ (.A1(_18402_),
    .A2(_18423_),
    .B1_N(_18422_),
    .Y(_18747_));
 sky130_fd_sc_hd__nor3_2 _28506_ (.A(_16271_),
    .B(_17627_),
    .C(_18358_),
    .Y(_18748_));
 sky130_fd_sc_hd__buf_1 _28507_ (.A(_14388_),
    .X(_18749_));
 sky130_fd_sc_hd__a22o_2 _28508_ (.A1(_14628_),
    .A2(_17630_),
    .B1(_18101_),
    .B2(_18749_),
    .X(_18750_));
 sky130_fd_sc_hd__and2b_2 _28509_ (.A_N(_18748_),
    .B(_18750_),
    .X(_18751_));
 sky130_fd_sc_hd__nor2_2 _28510_ (.A(_16625_),
    .B(_18114_),
    .Y(_18752_));
 sky130_fd_sc_hd__xnor2_2 _28511_ (.A(_18751_),
    .B(_18752_),
    .Y(_18753_));
 sky130_fd_sc_hd__buf_1 _28512_ (.A(_15624_),
    .X(_18754_));
 sky130_fd_sc_hd__or3b_2 _28513_ (.A(_14357_),
    .B(_16616_),
    .C_N(_18364_),
    .X(_18756_));
 sky130_fd_sc_hd__nor2_2 _28514_ (.A(_14357_),
    .B(_16255_),
    .Y(_18757_));
 sky130_fd_sc_hd__a21o_2 _28515_ (.A1(_16268_),
    .A2(_16613_),
    .B1(_18757_),
    .X(_18758_));
 sky130_fd_sc_hd__nand4_2 _28516_ (.A(_18754_),
    .B(_17393_),
    .C(_18756_),
    .D(_18758_),
    .Y(_18759_));
 sky130_fd_sc_hd__a22o_2 _28517_ (.A1(_18754_),
    .A2(_17393_),
    .B1(_18756_),
    .B2(_18758_),
    .X(_18760_));
 sky130_fd_sc_hd__a31o_2 _28518_ (.A1(_14629_),
    .A2(_17394_),
    .A3(_18366_),
    .B1(_18365_),
    .X(_18761_));
 sky130_fd_sc_hd__and3_2 _28519_ (.A(_18759_),
    .B(_18760_),
    .C(_18761_),
    .X(_18762_));
 sky130_fd_sc_hd__a21oi_2 _28520_ (.A1(_18759_),
    .A2(_18760_),
    .B1(_18761_),
    .Y(_18763_));
 sky130_fd_sc_hd__nor2_2 _28521_ (.A(_18762_),
    .B(_18763_),
    .Y(_18764_));
 sky130_fd_sc_hd__xnor2_2 _28522_ (.A(_18753_),
    .B(_18764_),
    .Y(_18765_));
 sky130_fd_sc_hd__nand2_2 _28523_ (.A(_18381_),
    .B(_18385_),
    .Y(_18767_));
 sky130_fd_sc_hd__a21bo_2 _28524_ (.A1(_18407_),
    .A2(_18409_),
    .B1_N(_18406_),
    .X(_18768_));
 sky130_fd_sc_hd__nor2_2 _28525_ (.A(_15211_),
    .B(_16237_),
    .Y(_18769_));
 sky130_fd_sc_hd__xnor2_2 _28526_ (.A(_18380_),
    .B(_18769_),
    .Y(_18770_));
 sky130_fd_sc_hd__nor2_2 _28527_ (.A(_14352_),
    .B(_15834_),
    .Y(_18771_));
 sky130_fd_sc_hd__xnor2_2 _28528_ (.A(_18770_),
    .B(_18771_),
    .Y(_18772_));
 sky130_fd_sc_hd__xor2_2 _28529_ (.A(_18768_),
    .B(_18772_),
    .X(_18773_));
 sky130_fd_sc_hd__xor2_2 _28530_ (.A(_18767_),
    .B(_18773_),
    .X(_18774_));
 sky130_fd_sc_hd__and2_2 _28531_ (.A(_18387_),
    .B(_18389_),
    .X(_18775_));
 sky130_fd_sc_hd__xnor2_2 _28532_ (.A(_18774_),
    .B(_18775_),
    .Y(_18776_));
 sky130_fd_sc_hd__xnor2_2 _28533_ (.A(_18765_),
    .B(_18776_),
    .Y(_18778_));
 sky130_fd_sc_hd__xnor2_2 _28534_ (.A(_18747_),
    .B(_18778_),
    .Y(_18779_));
 sky130_fd_sc_hd__xnor2_2 _28535_ (.A(_18746_),
    .B(_18779_),
    .Y(_18780_));
 sky130_fd_sc_hd__or2b_2 _28536_ (.A(_18418_),
    .B_N(_18420_),
    .X(_18781_));
 sky130_fd_sc_hd__or2b_2 _28537_ (.A(_18427_),
    .B_N(_18434_),
    .X(_18782_));
 sky130_fd_sc_hd__o21ai_2 _28538_ (.A1(_18428_),
    .A2(_18433_),
    .B1(_18782_),
    .Y(_18783_));
 sky130_fd_sc_hd__nor2_2 _28539_ (.A(_15168_),
    .B(_15004_),
    .Y(_18784_));
 sky130_fd_sc_hd__and3_2 _28540_ (.A(_15208_),
    .B(_14608_),
    .C(_18784_),
    .X(_18785_));
 sky130_fd_sc_hd__a21oi_2 _28541_ (.A1(_15208_),
    .A2(_14608_),
    .B1(_18784_),
    .Y(_18786_));
 sky130_fd_sc_hd__nor2_2 _28542_ (.A(_18785_),
    .B(_18786_),
    .Y(_18787_));
 sky130_fd_sc_hd__nor2_2 _28543_ (.A(_15648_),
    .B(_14949_),
    .Y(_18789_));
 sky130_fd_sc_hd__xnor2_2 _28544_ (.A(_18787_),
    .B(_18789_),
    .Y(_18790_));
 sky130_fd_sc_hd__buf_1 _28545_ (.A(_14612_),
    .X(_18791_));
 sky130_fd_sc_hd__nand2_2 _28546_ (.A(_13887_),
    .B(_15672_),
    .Y(_18792_));
 sky130_fd_sc_hd__a32o_2 _28547_ (.A1(_13888_),
    .A2(_15224_),
    .A3(_15226_),
    .B1(_15672_),
    .B2(_13543_),
    .X(_18793_));
 sky130_fd_sc_hd__o31ai_2 _28548_ (.A1(_18791_),
    .A2(_18181_),
    .A3(_18792_),
    .B1(_18793_),
    .Y(_18794_));
 sky130_fd_sc_hd__nand2_2 _28549_ (.A(_14392_),
    .B(_15679_),
    .Y(_18795_));
 sky130_fd_sc_hd__xnor2_2 _28550_ (.A(_18794_),
    .B(_18795_),
    .Y(_18796_));
 sky130_fd_sc_hd__and2_2 _28551_ (.A(_18412_),
    .B(_18414_),
    .X(_18797_));
 sky130_fd_sc_hd__xnor2_2 _28552_ (.A(_18796_),
    .B(_18797_),
    .Y(_18798_));
 sky130_fd_sc_hd__xor2_2 _28553_ (.A(_18790_),
    .B(_18798_),
    .X(_18799_));
 sky130_fd_sc_hd__xor2_2 _28554_ (.A(_18783_),
    .B(_18799_),
    .X(_18800_));
 sky130_fd_sc_hd__xnor2_2 _28555_ (.A(_18781_),
    .B(_18800_),
    .Y(_18801_));
 sky130_fd_sc_hd__a21bo_2 _28556_ (.A1(_18430_),
    .A2(_18432_),
    .B1_N(_18429_),
    .X(_18802_));
 sky130_fd_sc_hd__a31o_2 _28557_ (.A1(_15887_),
    .A2(_17488_),
    .A3(_18441_),
    .B1(_18438_),
    .X(_18803_));
 sky130_fd_sc_hd__or4_2 _28558_ (.A(_12848_),
    .B(_12850_),
    .C(_16988_),
    .D(_17007_),
    .X(_18804_));
 sky130_fd_sc_hd__a22o_2 _28559_ (.A1(_12846_),
    .A2(_17006_),
    .B1(_16680_),
    .B2(_14636_),
    .X(_18805_));
 sky130_fd_sc_hd__nand2_2 _28560_ (.A(_18804_),
    .B(_18805_),
    .Y(_18806_));
 sky130_fd_sc_hd__nor2_2 _28561_ (.A(_14625_),
    .B(_17696_),
    .Y(_18807_));
 sky130_fd_sc_hd__xnor2_2 _28562_ (.A(_18806_),
    .B(_18807_),
    .Y(_18808_));
 sky130_fd_sc_hd__xor2_2 _28563_ (.A(_18803_),
    .B(_18808_),
    .X(_18810_));
 sky130_fd_sc_hd__xnor2_2 _28564_ (.A(_18802_),
    .B(_18810_),
    .Y(_18811_));
 sky130_fd_sc_hd__nand2_2 _28565_ (.A(_15887_),
    .B(_17702_),
    .Y(_18812_));
 sky130_fd_sc_hd__and3_2 _28566_ (.A(_12243_),
    .B(_18205_),
    .C(_18439_),
    .X(_18813_));
 sky130_fd_sc_hd__a22o_2 _28567_ (.A1(_12243_),
    .A2(_17485_),
    .B1(_18205_),
    .B2(_14649_),
    .X(_18814_));
 sky130_fd_sc_hd__and2b_2 _28568_ (.A_N(_18813_),
    .B(_18814_),
    .X(_18815_));
 sky130_fd_sc_hd__xnor2_2 _28569_ (.A(_18812_),
    .B(_18815_),
    .Y(_18816_));
 sky130_fd_sc_hd__nor2_2 _28570_ (.A(_11793_),
    .B(_18211_),
    .Y(_18817_));
 sky130_fd_sc_hd__nor2_2 _28571_ (.A(iX[25]),
    .B(iX[57]),
    .Y(_18818_));
 sky130_fd_sc_hd__nand2_2 _28572_ (.A(iX[25]),
    .B(iX[57]),
    .Y(_18819_));
 sky130_fd_sc_hd__or2b_2 _28573_ (.A(_18818_),
    .B_N(_18819_),
    .X(_18821_));
 sky130_fd_sc_hd__and3_2 _28574_ (.A(_18451_),
    .B(_18454_),
    .C(_18821_),
    .X(_18822_));
 sky130_fd_sc_hd__a21oi_2 _28575_ (.A1(_18451_),
    .A2(_18454_),
    .B1(_18821_),
    .Y(_18823_));
 sky130_fd_sc_hd__or3_2 _28576_ (.A(_11566_),
    .B(_18822_),
    .C(_18823_),
    .X(_18824_));
 sky130_fd_sc_hd__xor2_2 _28577_ (.A(_18457_),
    .B(_18824_),
    .X(_18825_));
 sky130_fd_sc_hd__xnor2_2 _28578_ (.A(_18817_),
    .B(_18825_),
    .Y(_18826_));
 sky130_fd_sc_hd__a31o_2 _28579_ (.A1(_15675_),
    .A2(_18463_),
    .A3(_18461_),
    .B1(_18458_),
    .X(_18827_));
 sky130_fd_sc_hd__xor2_2 _28580_ (.A(_18826_),
    .B(_18827_),
    .X(_18828_));
 sky130_fd_sc_hd__xnor2_2 _28581_ (.A(_18816_),
    .B(_18828_),
    .Y(_18829_));
 sky130_fd_sc_hd__a21bo_2 _28582_ (.A1(_18442_),
    .A2(_18468_),
    .B1_N(_18467_),
    .X(_18830_));
 sky130_fd_sc_hd__xnor2_2 _28583_ (.A(_18829_),
    .B(_18830_),
    .Y(_18832_));
 sky130_fd_sc_hd__xnor2_2 _28584_ (.A(_18811_),
    .B(_18832_),
    .Y(_18833_));
 sky130_fd_sc_hd__a21bo_2 _28585_ (.A1(_18435_),
    .A2(_18474_),
    .B1_N(_18473_),
    .X(_18834_));
 sky130_fd_sc_hd__xor2_2 _28586_ (.A(_18833_),
    .B(_18834_),
    .X(_18835_));
 sky130_fd_sc_hd__xnor2_2 _28587_ (.A(_18801_),
    .B(_18835_),
    .Y(_18836_));
 sky130_fd_sc_hd__a21boi_2 _28588_ (.A1(_18425_),
    .A2(_18478_),
    .B1_N(_18477_),
    .Y(_18837_));
 sky130_fd_sc_hd__xnor2_2 _28589_ (.A(_18836_),
    .B(_18837_),
    .Y(_18838_));
 sky130_fd_sc_hd__xnor2_2 _28590_ (.A(_18780_),
    .B(_18838_),
    .Y(_18839_));
 sky130_fd_sc_hd__a21bo_2 _28591_ (.A1(_18400_),
    .A2(_18483_),
    .B1_N(_18482_),
    .X(_18840_));
 sky130_fd_sc_hd__xor2_2 _28592_ (.A(_18839_),
    .B(_18840_),
    .X(_18841_));
 sky130_fd_sc_hd__xnor2_2 _28593_ (.A(_18745_),
    .B(_18841_),
    .Y(_18843_));
 sky130_fd_sc_hd__a21bo_2 _28594_ (.A1(_18354_),
    .A2(_18487_),
    .B1_N(_18486_),
    .X(_18844_));
 sky130_fd_sc_hd__xnor2_2 _28595_ (.A(_18843_),
    .B(_18844_),
    .Y(_18845_));
 sky130_fd_sc_hd__xor2_2 _28596_ (.A(_18352_),
    .B(_18845_),
    .X(_18846_));
 sky130_fd_sc_hd__a21boi_2 _28597_ (.A1(_18322_),
    .A2(_18491_),
    .B1_N(_18490_),
    .Y(_18847_));
 sky130_fd_sc_hd__xor2_2 _28598_ (.A(_18846_),
    .B(_18847_),
    .X(_18848_));
 sky130_fd_sc_hd__nor2_2 _28599_ (.A(_18495_),
    .B(_18848_),
    .Y(_18849_));
 sky130_fd_sc_hd__and2_2 _28600_ (.A(_18495_),
    .B(_18848_),
    .X(_18850_));
 sky130_fd_sc_hd__nor2_2 _28601_ (.A(_18849_),
    .B(_18850_),
    .Y(_18851_));
 sky130_fd_sc_hd__nand3_2 _28602_ (.A(_18715_),
    .B(_18716_),
    .C(_18851_),
    .Y(_18852_));
 sky130_fd_sc_hd__a21o_2 _28603_ (.A1(_18715_),
    .A2(_18716_),
    .B1(_18851_),
    .X(_18854_));
 sky130_fd_sc_hd__and2_2 _28604_ (.A(_18640_),
    .B(_18641_),
    .X(_18855_));
 sky130_fd_sc_hd__nor2_2 _28605_ (.A(_18637_),
    .B(_18638_),
    .Y(_18856_));
 sky130_fd_sc_hd__nor2_2 _28606_ (.A(_18510_),
    .B(_18639_),
    .Y(_18857_));
 sky130_fd_sc_hd__a21oi_2 _28607_ (.A1(_18513_),
    .A2(_18515_),
    .B1(_18529_),
    .Y(_18858_));
 sky130_fd_sc_hd__or2b_2 _28608_ (.A(_18521_),
    .B_N(_18520_),
    .X(_18859_));
 sky130_fd_sc_hd__nand2_2 _28609_ (.A(_18522_),
    .B(_18528_),
    .Y(_18860_));
 sky130_fd_sc_hd__and4_2 _28610_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[54]),
    .D(iX[55]),
    .X(_18861_));
 sky130_fd_sc_hd__a22oi_2 _28611_ (.A1(iY[35]),
    .A2(iX[54]),
    .B1(iX[55]),
    .B2(iY[34]),
    .Y(_18862_));
 sky130_fd_sc_hd__nor2_2 _28612_ (.A(_18861_),
    .B(_18862_),
    .Y(_18863_));
 sky130_fd_sc_hd__nand2_2 _28613_ (.A(iY[33]),
    .B(iX[56]),
    .Y(_18865_));
 sky130_fd_sc_hd__xnor2_2 _28614_ (.A(_18863_),
    .B(_18865_),
    .Y(_18866_));
 sky130_fd_sc_hd__o21ba_2 _28615_ (.A1(_18517_),
    .A2(_18519_),
    .B1_N(_18516_),
    .X(_18867_));
 sky130_fd_sc_hd__xnor2_2 _28616_ (.A(_18866_),
    .B(_18867_),
    .Y(_18868_));
 sky130_fd_sc_hd__and4_2 _28617_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[53]),
    .D(iX[57]),
    .X(_18869_));
 sky130_fd_sc_hd__a22oi_2 _28618_ (.A1(iY[36]),
    .A2(iX[53]),
    .B1(iX[57]),
    .B2(iY[32]),
    .Y(_18870_));
 sky130_fd_sc_hd__nor2_2 _28619_ (.A(_18869_),
    .B(_18870_),
    .Y(_18871_));
 sky130_fd_sc_hd__nand2_2 _28620_ (.A(iY[37]),
    .B(iX[52]),
    .Y(_18872_));
 sky130_fd_sc_hd__xnor2_2 _28621_ (.A(_18871_),
    .B(_18872_),
    .Y(_18873_));
 sky130_fd_sc_hd__nand2_2 _28622_ (.A(_18868_),
    .B(_18873_),
    .Y(_18874_));
 sky130_fd_sc_hd__or2_2 _28623_ (.A(_18868_),
    .B(_18873_),
    .X(_18876_));
 sky130_fd_sc_hd__nand2_2 _28624_ (.A(_18874_),
    .B(_18876_),
    .Y(_18877_));
 sky130_fd_sc_hd__a21o_2 _28625_ (.A1(_18859_),
    .A2(_18860_),
    .B1(_18877_),
    .X(_18878_));
 sky130_fd_sc_hd__nand3_2 _28626_ (.A(_18859_),
    .B(_18860_),
    .C(_18877_),
    .Y(_18879_));
 sky130_fd_sc_hd__o21ba_2 _28627_ (.A1(_18535_),
    .A2(_18538_),
    .B1_N(_18534_),
    .X(_18880_));
 sky130_fd_sc_hd__o21ba_2 _28628_ (.A1(_18524_),
    .A2(_18527_),
    .B1_N(_18523_),
    .X(_18881_));
 sky130_fd_sc_hd__and4_2 _28629_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[50]),
    .D(iX[51]),
    .X(_18882_));
 sky130_fd_sc_hd__a22oi_2 _28630_ (.A1(iY[39]),
    .A2(iX[50]),
    .B1(iX[51]),
    .B2(iY[38]),
    .Y(_18883_));
 sky130_fd_sc_hd__nor2_2 _28631_ (.A(_18882_),
    .B(_18883_),
    .Y(_18884_));
 sky130_fd_sc_hd__nand2_2 _28632_ (.A(iY[40]),
    .B(iX[49]),
    .Y(_18885_));
 sky130_fd_sc_hd__xnor2_2 _28633_ (.A(_18884_),
    .B(_18885_),
    .Y(_18887_));
 sky130_fd_sc_hd__xnor2_2 _28634_ (.A(_18881_),
    .B(_18887_),
    .Y(_18888_));
 sky130_fd_sc_hd__xnor2_2 _28635_ (.A(_18880_),
    .B(_18888_),
    .Y(_18889_));
 sky130_fd_sc_hd__nand3_2 _28636_ (.A(_18878_),
    .B(_18879_),
    .C(_18889_),
    .Y(_18890_));
 sky130_fd_sc_hd__a21o_2 _28637_ (.A1(_18878_),
    .A2(_18879_),
    .B1(_18889_),
    .X(_18891_));
 sky130_fd_sc_hd__o211a_2 _28638_ (.A1(_18858_),
    .A2(_18542_),
    .B1(_18890_),
    .C1(_18891_),
    .X(_18892_));
 sky130_fd_sc_hd__a211oi_2 _28639_ (.A1(_18890_),
    .A2(_18891_),
    .B1(_18858_),
    .C1(_18542_),
    .Y(_18893_));
 sky130_fd_sc_hd__or2_2 _28640_ (.A(_18892_),
    .B(_18893_),
    .X(_18894_));
 sky130_fd_sc_hd__and2b_2 _28641_ (.A_N(_18562_),
    .B(_18561_),
    .X(_18895_));
 sky130_fd_sc_hd__a21o_2 _28642_ (.A1(_18555_),
    .A2(_18563_),
    .B1(_18895_),
    .X(_18896_));
 sky130_fd_sc_hd__or2b_2 _28643_ (.A(_18533_),
    .B_N(_18539_),
    .X(_18898_));
 sky130_fd_sc_hd__or2b_2 _28644_ (.A(_18532_),
    .B_N(_18540_),
    .X(_18899_));
 sky130_fd_sc_hd__and4_2 _28645_ (.A(iX[44]),
    .B(iY[44]),
    .C(iX[45]),
    .D(iY[45]),
    .X(_18900_));
 sky130_fd_sc_hd__a22oi_2 _28646_ (.A1(iY[44]),
    .A2(iX[45]),
    .B1(iY[45]),
    .B2(iX[44]),
    .Y(_18901_));
 sky130_fd_sc_hd__nor2_2 _28647_ (.A(_18900_),
    .B(_18901_),
    .Y(_18902_));
 sky130_fd_sc_hd__nand2_2 _28648_ (.A(iX[43]),
    .B(iY[46]),
    .Y(_18903_));
 sky130_fd_sc_hd__xnor2_2 _28649_ (.A(_18902_),
    .B(_18903_),
    .Y(_18904_));
 sky130_fd_sc_hd__and4_2 _28650_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[47]),
    .D(iX[48]),
    .X(_18905_));
 sky130_fd_sc_hd__a22oi_2 _28651_ (.A1(iY[42]),
    .A2(iX[47]),
    .B1(iX[48]),
    .B2(iY[41]),
    .Y(_18906_));
 sky130_fd_sc_hd__and4bb_2 _28652_ (.A_N(_18905_),
    .B_N(_18906_),
    .C(iY[43]),
    .D(iX[46]),
    .X(_18907_));
 sky130_fd_sc_hd__o2bb2a_2 _28653_ (.A1_N(iY[43]),
    .A2_N(iX[46]),
    .B1(_18905_),
    .B2(_18906_),
    .X(_18909_));
 sky130_fd_sc_hd__nor2_2 _28654_ (.A(_18907_),
    .B(_18909_),
    .Y(_18910_));
 sky130_fd_sc_hd__o21ba_2 _28655_ (.A1(_18557_),
    .A2(_18560_),
    .B1_N(_18556_),
    .X(_18911_));
 sky130_fd_sc_hd__xnor2_2 _28656_ (.A(_18910_),
    .B(_18911_),
    .Y(_18912_));
 sky130_fd_sc_hd__and2_2 _28657_ (.A(_18904_),
    .B(_18912_),
    .X(_18913_));
 sky130_fd_sc_hd__nor2_2 _28658_ (.A(_18904_),
    .B(_18912_),
    .Y(_18914_));
 sky130_fd_sc_hd__or2_2 _28659_ (.A(_18913_),
    .B(_18914_),
    .X(_18915_));
 sky130_fd_sc_hd__a21o_2 _28660_ (.A1(_18898_),
    .A2(_18899_),
    .B1(_18915_),
    .X(_18916_));
 sky130_fd_sc_hd__nand3_2 _28661_ (.A(_18898_),
    .B(_18899_),
    .C(_18915_),
    .Y(_18917_));
 sky130_fd_sc_hd__nand3_2 _28662_ (.A(_18896_),
    .B(_18916_),
    .C(_18917_),
    .Y(_18918_));
 sky130_fd_sc_hd__a21o_2 _28663_ (.A1(_18916_),
    .A2(_18917_),
    .B1(_18896_),
    .X(_18920_));
 sky130_fd_sc_hd__nand2_2 _28664_ (.A(_18918_),
    .B(_18920_),
    .Y(_18921_));
 sky130_fd_sc_hd__xor2_2 _28665_ (.A(_18894_),
    .B(_18921_),
    .X(_18922_));
 sky130_fd_sc_hd__a21bo_2 _28666_ (.A1(_18544_),
    .A2(_18545_),
    .B1_N(_18571_),
    .X(_18923_));
 sky130_fd_sc_hd__xnor2_2 _28667_ (.A(_18922_),
    .B(_18923_),
    .Y(_18924_));
 sky130_fd_sc_hd__and4_2 _28668_ (.A(iX[35]),
    .B(iX[36]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_18925_));
 sky130_fd_sc_hd__a22oi_2 _28669_ (.A1(iX[36]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[35]),
    .Y(_18926_));
 sky130_fd_sc_hd__nor2_2 _28670_ (.A(_18925_),
    .B(_18926_),
    .Y(_18927_));
 sky130_fd_sc_hd__nand2_2 _28671_ (.A(iX[34]),
    .B(iY[55]),
    .Y(_18928_));
 sky130_fd_sc_hd__xnor2_2 _28672_ (.A(_18927_),
    .B(_18928_),
    .Y(_18929_));
 sky130_fd_sc_hd__and4_2 _28673_ (.A(iX[38]),
    .B(iX[39]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_00001_));
 sky130_fd_sc_hd__a22oi_2 _28674_ (.A1(iX[39]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[38]),
    .Y(_00002_));
 sky130_fd_sc_hd__nor2_2 _28675_ (.A(_00001_),
    .B(_00002_),
    .Y(_00003_));
 sky130_fd_sc_hd__nand2_2 _28676_ (.A(iX[37]),
    .B(iY[52]),
    .Y(_00004_));
 sky130_fd_sc_hd__xnor2_2 _28677_ (.A(_00003_),
    .B(_00004_),
    .Y(_00005_));
 sky130_fd_sc_hd__o21ba_2 _28678_ (.A1(_18584_),
    .A2(_18586_),
    .B1_N(_18583_),
    .X(_00006_));
 sky130_fd_sc_hd__xnor2_2 _28679_ (.A(_00005_),
    .B(_00006_),
    .Y(_00007_));
 sky130_fd_sc_hd__nand2_2 _28680_ (.A(_18929_),
    .B(_00007_),
    .Y(_00008_));
 sky130_fd_sc_hd__or2_2 _28681_ (.A(_18929_),
    .B(_00007_),
    .X(_00009_));
 sky130_fd_sc_hd__nand2_2 _28682_ (.A(_00008_),
    .B(_00009_),
    .Y(_00010_));
 sky130_fd_sc_hd__or3_2 _28683_ (.A(_18596_),
    .B(_18599_),
    .C(_18600_),
    .X(_00012_));
 sky130_fd_sc_hd__o21ba_2 _28684_ (.A1(_18552_),
    .A2(_18554_),
    .B1_N(_18551_),
    .X(_00013_));
 sky130_fd_sc_hd__and4_2 _28685_ (.A(iX[41]),
    .B(iX[42]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_00014_));
 sky130_fd_sc_hd__a22oi_2 _28686_ (.A1(iX[42]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[41]),
    .Y(_00015_));
 sky130_fd_sc_hd__and4bb_2 _28687_ (.A_N(_00014_),
    .B_N(_00015_),
    .C(iX[40]),
    .D(iY[49]),
    .X(_00016_));
 sky130_fd_sc_hd__o2bb2a_2 _28688_ (.A1_N(iX[40]),
    .A2_N(iY[49]),
    .B1(_00014_),
    .B2(_00015_),
    .X(_00017_));
 sky130_fd_sc_hd__nor2_2 _28689_ (.A(_00016_),
    .B(_00017_),
    .Y(_00018_));
 sky130_fd_sc_hd__xnor2_2 _28690_ (.A(_00013_),
    .B(_00018_),
    .Y(_00019_));
 sky130_fd_sc_hd__o21ai_2 _28691_ (.A1(_18597_),
    .A2(_18599_),
    .B1(_00019_),
    .Y(_00020_));
 sky130_fd_sc_hd__or3_2 _28692_ (.A(_18597_),
    .B(_18599_),
    .C(_00019_),
    .X(_00021_));
 sky130_fd_sc_hd__nand2_2 _28693_ (.A(_00020_),
    .B(_00021_),
    .Y(_00023_));
 sky130_fd_sc_hd__a21oi_2 _28694_ (.A1(_00012_),
    .A2(_18604_),
    .B1(_00023_),
    .Y(_00024_));
 sky130_fd_sc_hd__and3_2 _28695_ (.A(_00012_),
    .B(_18604_),
    .C(_00023_),
    .X(_00025_));
 sky130_fd_sc_hd__or3_2 _28696_ (.A(_00010_),
    .B(_00024_),
    .C(_00025_),
    .X(_00026_));
 sky130_fd_sc_hd__o21ai_2 _28697_ (.A1(_00024_),
    .A2(_00025_),
    .B1(_00010_),
    .Y(_00027_));
 sky130_fd_sc_hd__o211a_2 _28698_ (.A1(_18565_),
    .A2(_18568_),
    .B1(_00026_),
    .C1(_00027_),
    .X(_00028_));
 sky130_fd_sc_hd__inv_2 _28699_ (.A(_00028_),
    .Y(_00029_));
 sky130_fd_sc_hd__a211o_2 _28700_ (.A1(_00026_),
    .A2(_00027_),
    .B1(_18565_),
    .C1(_18568_),
    .X(_00030_));
 sky130_fd_sc_hd__o211a_2 _28701_ (.A1(_18607_),
    .A2(_18609_),
    .B1(_00029_),
    .C1(_00030_),
    .X(_00031_));
 sky130_fd_sc_hd__a211oi_2 _28702_ (.A1(_00029_),
    .A2(_00030_),
    .B1(_18607_),
    .C1(_18609_),
    .Y(_00032_));
 sky130_fd_sc_hd__nor2_2 _28703_ (.A(_00031_),
    .B(_00032_),
    .Y(_00034_));
 sky130_fd_sc_hd__xnor2_2 _28704_ (.A(_18924_),
    .B(_00034_),
    .Y(_00035_));
 sky130_fd_sc_hd__o21a_2 _28705_ (.A1(_18574_),
    .A2(_18616_),
    .B1(_00035_),
    .X(_00036_));
 sky130_fd_sc_hd__nor3_2 _28706_ (.A(_18574_),
    .B(_18616_),
    .C(_00035_),
    .Y(_00037_));
 sky130_fd_sc_hd__and3_2 _28707_ (.A(_17816_),
    .B(_18061_),
    .C(_18629_),
    .X(_00038_));
 sky130_fd_sc_hd__and2_2 _28708_ (.A(_18587_),
    .B(_18588_),
    .X(_00039_));
 sky130_fd_sc_hd__a31o_2 _28709_ (.A1(iX[33]),
    .A2(iY[55]),
    .A3(_18579_),
    .B1(_18577_),
    .X(_00040_));
 sky130_fd_sc_hd__a22o_2 _28710_ (.A1(iX[33]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[32]),
    .X(_00041_));
 sky130_fd_sc_hd__and4_2 _28711_ (.A(iX[33]),
    .B(iX[32]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_00042_));
 sky130_fd_sc_hd__inv_2 _28712_ (.A(_00042_),
    .Y(_00043_));
 sky130_fd_sc_hd__and3_2 _28713_ (.A(_00040_),
    .B(_00041_),
    .C(_00043_),
    .X(_00045_));
 sky130_fd_sc_hd__a21oi_2 _28714_ (.A1(_00041_),
    .A2(_00043_),
    .B1(_00040_),
    .Y(_00046_));
 sky130_fd_sc_hd__nor2_2 _28715_ (.A(_00045_),
    .B(_00046_),
    .Y(_00047_));
 sky130_fd_sc_hd__o21ai_2 _28716_ (.A1(_00039_),
    .A2(_18590_),
    .B1(_00047_),
    .Y(_00048_));
 sky130_fd_sc_hd__or3_2 _28717_ (.A(_00039_),
    .B(_18590_),
    .C(_00047_),
    .X(_00049_));
 sky130_fd_sc_hd__and2_2 _28718_ (.A(_00048_),
    .B(_00049_),
    .X(_00050_));
 sky130_fd_sc_hd__nand2_2 _28719_ (.A(_18623_),
    .B(_00050_),
    .Y(_00051_));
 sky130_fd_sc_hd__or2_2 _28720_ (.A(_18623_),
    .B(_00050_),
    .X(_00052_));
 sky130_fd_sc_hd__nand2_2 _28721_ (.A(_00051_),
    .B(_00052_),
    .Y(_00053_));
 sky130_fd_sc_hd__nor2_2 _28722_ (.A(_18627_),
    .B(_00053_),
    .Y(_00054_));
 sky130_fd_sc_hd__and2_2 _28723_ (.A(_18627_),
    .B(_00053_),
    .X(_00056_));
 sky130_fd_sc_hd__nor2_2 _28724_ (.A(_00054_),
    .B(_00056_),
    .Y(_00057_));
 sky130_fd_sc_hd__o21a_2 _28725_ (.A1(_18611_),
    .A2(_18614_),
    .B1(_00057_),
    .X(_00058_));
 sky130_fd_sc_hd__nor3_2 _28726_ (.A(_18611_),
    .B(_18614_),
    .C(_00057_),
    .Y(_00059_));
 sky130_fd_sc_hd__nor2_2 _28727_ (.A(_00058_),
    .B(_00059_),
    .Y(_00060_));
 sky130_fd_sc_hd__xnor2_2 _28728_ (.A(_00038_),
    .B(_00060_),
    .Y(_00061_));
 sky130_fd_sc_hd__nor3_2 _28729_ (.A(_00036_),
    .B(_00037_),
    .C(_00061_),
    .Y(_00062_));
 sky130_fd_sc_hd__o21a_2 _28730_ (.A1(_00036_),
    .A2(_00037_),
    .B1(_00061_),
    .X(_00063_));
 sky130_fd_sc_hd__nor2_2 _28731_ (.A(_00062_),
    .B(_00063_),
    .Y(_00064_));
 sky130_fd_sc_hd__o21ai_2 _28732_ (.A1(_18618_),
    .A2(_18634_),
    .B1(_00064_),
    .Y(_00065_));
 sky130_fd_sc_hd__or3_2 _28733_ (.A(_18618_),
    .B(_18634_),
    .C(_00064_),
    .X(_00067_));
 sky130_fd_sc_hd__nand3_2 _28734_ (.A(_18631_),
    .B(_00065_),
    .C(_00067_),
    .Y(_00068_));
 sky130_fd_sc_hd__a21o_2 _28735_ (.A1(_00065_),
    .A2(_00067_),
    .B1(_18631_),
    .X(_00069_));
 sky130_fd_sc_hd__o211ai_2 _28736_ (.A1(_18856_),
    .A2(_18857_),
    .B1(_00068_),
    .C1(_00069_),
    .Y(_00070_));
 sky130_fd_sc_hd__a211o_2 _28737_ (.A1(_00068_),
    .A2(_00069_),
    .B1(_18856_),
    .C1(_18857_),
    .X(_00071_));
 sky130_fd_sc_hd__and3_2 _28738_ (.A(_18855_),
    .B(_00070_),
    .C(_00071_),
    .X(_00072_));
 sky130_fd_sc_hd__a21oi_2 _28739_ (.A1(_00070_),
    .A2(_00071_),
    .B1(_18855_),
    .Y(_00073_));
 sky130_fd_sc_hd__nor2_2 _28740_ (.A(_00072_),
    .B(_00073_),
    .Y(_00074_));
 sky130_fd_sc_hd__a21oi_2 _28741_ (.A1(_18508_),
    .A2(_18645_),
    .B1(_18643_),
    .Y(_00075_));
 sky130_fd_sc_hd__xnor2_2 _28742_ (.A(_00074_),
    .B(_00075_),
    .Y(_00076_));
 sky130_fd_sc_hd__and3_2 _28743_ (.A(_18852_),
    .B(_18854_),
    .C(_00076_),
    .X(_00078_));
 sky130_fd_sc_hd__a21oi_2 _28744_ (.A1(_18852_),
    .A2(_18854_),
    .B1(_00076_),
    .Y(_00079_));
 sky130_fd_sc_hd__or3_2 _28745_ (.A(oO[25]),
    .B(_00078_),
    .C(_00079_),
    .X(_00080_));
 sky130_fd_sc_hd__o21ai_2 _28746_ (.A1(_00078_),
    .A2(_00079_),
    .B1(oO[25]),
    .Y(_00081_));
 sky130_fd_sc_hd__and2b_2 _28747_ (.A_N(_18647_),
    .B(_18500_),
    .X(_00082_));
 sky130_fd_sc_hd__a21o_2 _28748_ (.A1(_09530_),
    .A2(_18648_),
    .B1(_00082_),
    .X(_00083_));
 sky130_fd_sc_hd__and3_2 _28749_ (.A(_00080_),
    .B(_00081_),
    .C(_00083_),
    .X(_00084_));
 sky130_fd_sc_hd__a21oi_2 _28750_ (.A1(_00080_),
    .A2(_00081_),
    .B1(_00083_),
    .Y(_00085_));
 sky130_fd_sc_hd__or2_2 _28751_ (.A(_00084_),
    .B(_00085_),
    .X(_00086_));
 sky130_fd_sc_hd__or2_2 _28752_ (.A(_18649_),
    .B(_18651_),
    .X(_00087_));
 sky130_fd_sc_hd__o21a_2 _28753_ (.A1(_18652_),
    .A2(_18656_),
    .B1(_00087_),
    .X(_00089_));
 sky130_fd_sc_hd__xnor2_2 _28754_ (.A(_00086_),
    .B(_00089_),
    .Y(_00090_));
 sky130_fd_sc_hd__and2_2 _28755_ (.A(_18714_),
    .B(_00090_),
    .X(_00091_));
 sky130_fd_sc_hd__nor2_2 _28756_ (.A(_18714_),
    .B(_00090_),
    .Y(_00092_));
 sky130_fd_sc_hd__or2_2 _28757_ (.A(_00091_),
    .B(_00092_),
    .X(_00093_));
 sky130_fd_sc_hd__inv_2 _28758_ (.A(_00093_),
    .Y(_00094_));
 sky130_fd_sc_hd__and2b_2 _28759_ (.A_N(_18312_),
    .B(_18658_),
    .X(_00095_));
 sky130_fd_sc_hd__o21ba_2 _28760_ (.A1(_18659_),
    .A2(_18669_),
    .B1_N(_00095_),
    .X(_00096_));
 sky130_fd_sc_hd__xnor2_2 _28761_ (.A(_00094_),
    .B(_00096_),
    .Y(oO[57]));
 sky130_fd_sc_hd__o211a_2 _28762_ (.A1(_18665_),
    .A2(_18667_),
    .B1(_00094_),
    .C1(_18660_),
    .X(_00097_));
 sky130_fd_sc_hd__nor2_2 _28763_ (.A(_00095_),
    .B(_00092_),
    .Y(_00099_));
 sky130_fd_sc_hd__nor2_2 _28764_ (.A(_00091_),
    .B(_00099_),
    .Y(_00100_));
 sky130_fd_sc_hd__o221a_2 _28765_ (.A1(_18706_),
    .A2(_18707_),
    .B1(_18708_),
    .B2(_18670_),
    .C1(_18713_),
    .X(_00101_));
 sky130_fd_sc_hd__or2b_2 _28766_ (.A(_18677_),
    .B_N(_18676_),
    .X(_00102_));
 sky130_fd_sc_hd__nand2_2 _28767_ (.A(iY[28]),
    .B(iX[30]),
    .Y(_00103_));
 sky130_fd_sc_hd__nand2_2 _28768_ (.A(iY[27]),
    .B(iX[31]),
    .Y(_00104_));
 sky130_fd_sc_hd__and4_2 _28769_ (.A(iY[27]),
    .B(iY[28]),
    .C(iX[30]),
    .D(iX[31]),
    .X(_00105_));
 sky130_fd_sc_hd__a21o_2 _28770_ (.A1(_00103_),
    .A2(_00104_),
    .B1(_00105_),
    .X(_00106_));
 sky130_fd_sc_hd__nand2_2 _28771_ (.A(iX[29]),
    .B(iY[29]),
    .Y(_00107_));
 sky130_fd_sc_hd__xor2_2 _28772_ (.A(_00106_),
    .B(_00107_),
    .X(_00108_));
 sky130_fd_sc_hd__o21ba_2 _28773_ (.A1(_18673_),
    .A2(_18675_),
    .B1_N(_18672_),
    .X(_00110_));
 sky130_fd_sc_hd__xnor2_2 _28774_ (.A(_00108_),
    .B(_00110_),
    .Y(_00111_));
 sky130_fd_sc_hd__nand2_2 _28775_ (.A(iX[28]),
    .B(iY[30]),
    .Y(_00112_));
 sky130_fd_sc_hd__xor2_2 _28776_ (.A(_00111_),
    .B(_00112_),
    .X(_00113_));
 sky130_fd_sc_hd__a21oi_2 _28777_ (.A1(_00102_),
    .A2(_18680_),
    .B1(_00113_),
    .Y(_00114_));
 sky130_fd_sc_hd__and3_2 _28778_ (.A(_00102_),
    .B(_18680_),
    .C(_00113_),
    .X(_00115_));
 sky130_fd_sc_hd__nor2_2 _28779_ (.A(_00114_),
    .B(_00115_),
    .Y(_00116_));
 sky130_fd_sc_hd__nand2_2 _28780_ (.A(iX[27]),
    .B(iY[31]),
    .Y(_00117_));
 sky130_fd_sc_hd__xnor2_2 _28781_ (.A(_00116_),
    .B(_00117_),
    .Y(_00118_));
 sky130_fd_sc_hd__o211a_2 _28782_ (.A1(_17543_),
    .A2(_18296_),
    .B1(iY[26]),
    .C1(iX[31]),
    .X(_00119_));
 sky130_fd_sc_hd__nand2_2 _28783_ (.A(_00118_),
    .B(_00119_),
    .Y(_00121_));
 sky130_fd_sc_hd__or2_2 _28784_ (.A(_00118_),
    .B(_00119_),
    .X(_00122_));
 sky130_fd_sc_hd__and2_2 _28785_ (.A(_00121_),
    .B(_00122_),
    .X(_00123_));
 sky130_fd_sc_hd__a22o_2 _28786_ (.A1(_18691_),
    .A2(_18690_),
    .B1(_18693_),
    .B2(_18688_),
    .X(_00124_));
 sky130_fd_sc_hd__xor2_2 _28787_ (.A(_00123_),
    .B(_00124_),
    .X(_00125_));
 sky130_fd_sc_hd__a21o_2 _28788_ (.A1(_18302_),
    .A2(_18698_),
    .B1(_18696_),
    .X(_00126_));
 sky130_fd_sc_hd__xnor2_2 _28789_ (.A(_00125_),
    .B(_00126_),
    .Y(_00127_));
 sky130_fd_sc_hd__a21oi_2 _28790_ (.A1(_18683_),
    .A2(_18687_),
    .B1(_00127_),
    .Y(_00128_));
 sky130_fd_sc_hd__and3_2 _28791_ (.A(_18683_),
    .B(_18687_),
    .C(_00127_),
    .X(_00129_));
 sky130_fd_sc_hd__or2_2 _28792_ (.A(_00128_),
    .B(_00129_),
    .X(_00130_));
 sky130_fd_sc_hd__a21oi_2 _28793_ (.A1(_18699_),
    .A2(_18698_),
    .B1(_18703_),
    .Y(_00132_));
 sky130_fd_sc_hd__nor2_2 _28794_ (.A(_00130_),
    .B(_00132_),
    .Y(_00133_));
 sky130_fd_sc_hd__and2_2 _28795_ (.A(_00130_),
    .B(_00132_),
    .X(_00134_));
 sky130_fd_sc_hd__or2_2 _28796_ (.A(_00133_),
    .B(_00134_),
    .X(_00135_));
 sky130_fd_sc_hd__nor2_2 _28797_ (.A(_00101_),
    .B(_00135_),
    .Y(_00136_));
 sky130_fd_sc_hd__and2_2 _28798_ (.A(_00101_),
    .B(_00135_),
    .X(_00137_));
 sky130_fd_sc_hd__nor2_2 _28799_ (.A(_00136_),
    .B(_00137_),
    .Y(_00138_));
 sky130_fd_sc_hd__a21o_2 _28800_ (.A1(_18852_),
    .A2(_18854_),
    .B1(_00076_),
    .X(_00139_));
 sky130_fd_sc_hd__nor2_2 _28801_ (.A(_18846_),
    .B(_18847_),
    .Y(_00140_));
 sky130_fd_sc_hd__and2b_2 _28802_ (.A_N(_18843_),
    .B(_18844_),
    .X(_00141_));
 sky130_fd_sc_hd__and2b_2 _28803_ (.A_N(_18352_),
    .B(_18845_),
    .X(_00143_));
 sky130_fd_sc_hd__nor2_2 _28804_ (.A(_00141_),
    .B(_00143_),
    .Y(_00144_));
 sky130_fd_sc_hd__and2b_2 _28805_ (.A_N(_18717_),
    .B(_18742_),
    .X(_00145_));
 sky130_fd_sc_hd__a21oi_2 _28806_ (.A1(_18348_),
    .A2(_18743_),
    .B1(_00145_),
    .Y(_00146_));
 sky130_fd_sc_hd__or2_2 _28807_ (.A(_18718_),
    .B(_18741_),
    .X(_00147_));
 sky130_fd_sc_hd__and2b_2 _28808_ (.A_N(_18779_),
    .B(_18746_),
    .X(_00148_));
 sky130_fd_sc_hd__a21o_2 _28809_ (.A1(_18747_),
    .A2(_18778_),
    .B1(_00148_),
    .X(_00149_));
 sky130_fd_sc_hd__o21bai_2 _28810_ (.A1(_18753_),
    .A2(_18763_),
    .B1_N(_18762_),
    .Y(_00150_));
 sky130_fd_sc_hd__a31o_2 _28811_ (.A1(_15616_),
    .A2(_18326_),
    .A3(_18750_),
    .B1(_18748_),
    .X(_00151_));
 sky130_fd_sc_hd__or4b_2 _28812_ (.A(_11570_),
    .B(_16625_),
    .C(_18342_),
    .D_N(_18728_),
    .X(_00152_));
 sky130_fd_sc_hd__a22o_2 _28813_ (.A1(_15616_),
    .A2(_18732_),
    .B1(_18728_),
    .B2(_12838_),
    .X(_00154_));
 sky130_fd_sc_hd__nand2_2 _28814_ (.A(iY[26]),
    .B(iY[58]),
    .Y(_00155_));
 sky130_fd_sc_hd__or2_2 _28815_ (.A(iY[26]),
    .B(iY[58]),
    .X(_00156_));
 sky130_fd_sc_hd__nand2_2 _28816_ (.A(_00155_),
    .B(_00156_),
    .Y(_00157_));
 sky130_fd_sc_hd__a21oi_2 _28817_ (.A1(iY[24]),
    .A2(iY[56]),
    .B1(_18725_),
    .Y(_00158_));
 sky130_fd_sc_hd__o31a_2 _28818_ (.A1(_18333_),
    .A2(_18337_),
    .A3(_18339_),
    .B1(_00158_),
    .X(_00159_));
 sky130_fd_sc_hd__nor2_4 _28819_ (.A(_18724_),
    .B(_00159_),
    .Y(_00160_));
 sky130_fd_sc_hd__xnor2_2 _28820_ (.A(_00157_),
    .B(_00160_),
    .Y(_00161_));
 sky130_fd_sc_hd__buf_2 _28821_ (.A(_00161_),
    .X(_00162_));
 sky130_fd_sc_hd__nand4_2 _28822_ (.A(_14592_),
    .B(_00152_),
    .C(_00154_),
    .D(_00162_),
    .Y(_00163_));
 sky130_fd_sc_hd__a22o_2 _28823_ (.A1(_00152_),
    .A2(_00154_),
    .B1(_00161_),
    .B2(_14592_),
    .X(_00165_));
 sky130_fd_sc_hd__nand3_2 _28824_ (.A(_00151_),
    .B(_00163_),
    .C(_00165_),
    .Y(_00166_));
 sky130_fd_sc_hd__a21o_2 _28825_ (.A1(_00163_),
    .A2(_00165_),
    .B1(_00151_),
    .X(_00167_));
 sky130_fd_sc_hd__nand3_2 _28826_ (.A(_18735_),
    .B(_00166_),
    .C(_00167_),
    .Y(_00168_));
 sky130_fd_sc_hd__a21o_2 _28827_ (.A1(_00166_),
    .A2(_00167_),
    .B1(_18735_),
    .X(_00169_));
 sky130_fd_sc_hd__and3_2 _28828_ (.A(_00150_),
    .B(_00168_),
    .C(_00169_),
    .X(_00170_));
 sky130_fd_sc_hd__a21oi_2 _28829_ (.A1(_00168_),
    .A2(_00169_),
    .B1(_00150_),
    .Y(_00171_));
 sky130_fd_sc_hd__or2_2 _28830_ (.A(_00170_),
    .B(_00171_),
    .X(_00172_));
 sky130_fd_sc_hd__xor2_2 _28831_ (.A(_18737_),
    .B(_00172_),
    .X(_00173_));
 sky130_fd_sc_hd__a32oi_2 _28832_ (.A1(_18720_),
    .A2(_18737_),
    .A3(_18738_),
    .B1(_18740_),
    .B2(_18719_),
    .Y(_00174_));
 sky130_fd_sc_hd__xnor2_2 _28833_ (.A(_00173_),
    .B(_00174_),
    .Y(_00176_));
 sky130_fd_sc_hd__xor2_2 _28834_ (.A(_00149_),
    .B(_00176_),
    .X(_00177_));
 sky130_fd_sc_hd__xnor2_2 _28835_ (.A(_00147_),
    .B(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_2 _28836_ (.A(_18774_),
    .B(_18775_),
    .Y(_00179_));
 sky130_fd_sc_hd__or2_2 _28837_ (.A(_18774_),
    .B(_18775_),
    .X(_00180_));
 sky130_fd_sc_hd__a21bo_2 _28838_ (.A1(_18765_),
    .A2(_00179_),
    .B1_N(_00180_),
    .X(_00181_));
 sky130_fd_sc_hd__and2_2 _28839_ (.A(_18783_),
    .B(_18799_),
    .X(_00182_));
 sky130_fd_sc_hd__and2_2 _28840_ (.A(_18781_),
    .B(_18800_),
    .X(_00183_));
 sky130_fd_sc_hd__and4_2 _28841_ (.A(_14628_),
    .B(_15624_),
    .C(_17630_),
    .D(_18101_),
    .X(_00184_));
 sky130_fd_sc_hd__o22a_2 _28842_ (.A1(_18368_),
    .A2(_17408_),
    .B1(_17627_),
    .B2(_16271_),
    .X(_00185_));
 sky130_fd_sc_hd__or3_4 _28843_ (.A(_18120_),
    .B(_18110_),
    .C(_18112_),
    .X(_00187_));
 sky130_fd_sc_hd__o21a_2 _28844_ (.A1(_00184_),
    .A2(_00185_),
    .B1(_00187_),
    .X(_00188_));
 sky130_fd_sc_hd__or3_4 _28845_ (.A(_00184_),
    .B(_00185_),
    .C(_00187_),
    .X(_00189_));
 sky130_fd_sc_hd__nor2b_2 _28846_ (.A(_00188_),
    .B_N(_00189_),
    .Y(_00190_));
 sky130_fd_sc_hd__or3b_2 _28847_ (.A(_14352_),
    .B(_16617_),
    .C_N(_18757_),
    .X(_00191_));
 sky130_fd_sc_hd__nor2_2 _28848_ (.A(_14352_),
    .B(_16255_),
    .Y(_00192_));
 sky130_fd_sc_hd__a21o_2 _28849_ (.A1(_16277_),
    .A2(_16613_),
    .B1(_00192_),
    .X(_00193_));
 sky130_fd_sc_hd__nand2_2 _28850_ (.A(_00191_),
    .B(_00193_),
    .Y(_00194_));
 sky130_fd_sc_hd__buf_1 _28851_ (.A(_14343_),
    .X(_00195_));
 sky130_fd_sc_hd__or2_2 _28852_ (.A(_00195_),
    .B(_16922_),
    .X(_00196_));
 sky130_fd_sc_hd__xnor2_2 _28853_ (.A(_00194_),
    .B(_00196_),
    .Y(_00198_));
 sky130_fd_sc_hd__and2_2 _28854_ (.A(_18756_),
    .B(_18759_),
    .X(_00199_));
 sky130_fd_sc_hd__xor2_2 _28855_ (.A(_00198_),
    .B(_00199_),
    .X(_00200_));
 sky130_fd_sc_hd__xor2_2 _28856_ (.A(_00190_),
    .B(_00200_),
    .X(_00201_));
 sky130_fd_sc_hd__or2b_2 _28857_ (.A(_18772_),
    .B_N(_18768_),
    .X(_00202_));
 sky130_fd_sc_hd__or2b_2 _28858_ (.A(_18773_),
    .B_N(_18767_),
    .X(_00203_));
 sky130_fd_sc_hd__and2b_2 _28859_ (.A_N(_18380_),
    .B(_18769_),
    .X(_00204_));
 sky130_fd_sc_hd__a21o_2 _28860_ (.A1(_18770_),
    .A2(_18771_),
    .B1(_00204_),
    .X(_00205_));
 sky130_fd_sc_hd__a21o_2 _28861_ (.A1(_18787_),
    .A2(_18789_),
    .B1(_18785_),
    .X(_00206_));
 sky130_fd_sc_hd__nor2_2 _28862_ (.A(_15647_),
    .B(_15597_),
    .Y(_00207_));
 sky130_fd_sc_hd__o22a_2 _28863_ (.A1(_15647_),
    .A2(_16237_),
    .B1(_15598_),
    .B2(_15211_),
    .X(_00209_));
 sky130_fd_sc_hd__a21o_2 _28864_ (.A1(_18769_),
    .A2(_00207_),
    .B1(_00209_),
    .X(_00210_));
 sky130_fd_sc_hd__or2_2 _28865_ (.A(_14983_),
    .B(_15834_),
    .X(_00211_));
 sky130_fd_sc_hd__xor2_2 _28866_ (.A(_00210_),
    .B(_00211_),
    .X(_00212_));
 sky130_fd_sc_hd__xor2_2 _28867_ (.A(_00206_),
    .B(_00212_),
    .X(_00213_));
 sky130_fd_sc_hd__xnor2_2 _28868_ (.A(_00205_),
    .B(_00213_),
    .Y(_00214_));
 sky130_fd_sc_hd__a21o_2 _28869_ (.A1(_00202_),
    .A2(_00203_),
    .B1(_00214_),
    .X(_00215_));
 sky130_fd_sc_hd__nand3_2 _28870_ (.A(_00202_),
    .B(_00203_),
    .C(_00214_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand3_2 _28871_ (.A(_00201_),
    .B(_00215_),
    .C(_00216_),
    .Y(_00217_));
 sky130_fd_sc_hd__a21o_2 _28872_ (.A1(_00215_),
    .A2(_00216_),
    .B1(_00201_),
    .X(_00218_));
 sky130_fd_sc_hd__o211a_2 _28873_ (.A1(_00182_),
    .A2(_00183_),
    .B1(_00217_),
    .C1(_00218_),
    .X(_00220_));
 sky130_fd_sc_hd__a211oi_2 _28874_ (.A1(_00217_),
    .A2(_00218_),
    .B1(_00182_),
    .C1(_00183_),
    .Y(_00221_));
 sky130_fd_sc_hd__or2_2 _28875_ (.A(_00220_),
    .B(_00221_),
    .X(_00222_));
 sky130_fd_sc_hd__xnor2_2 _28876_ (.A(_00181_),
    .B(_00222_),
    .Y(_00223_));
 sky130_fd_sc_hd__or2_2 _28877_ (.A(_18790_),
    .B(_18798_),
    .X(_00224_));
 sky130_fd_sc_hd__o21a_2 _28878_ (.A1(_18796_),
    .A2(_18797_),
    .B1(_00224_),
    .X(_00225_));
 sky130_fd_sc_hd__and2_2 _28879_ (.A(_18803_),
    .B(_18808_),
    .X(_00226_));
 sky130_fd_sc_hd__and2_2 _28880_ (.A(_18802_),
    .B(_18810_),
    .X(_00227_));
 sky130_fd_sc_hd__nand2_2 _28881_ (.A(_14608_),
    .B(_16292_),
    .Y(_00228_));
 sky130_fd_sc_hd__nor2_2 _28882_ (.A(_15168_),
    .B(_14998_),
    .Y(_00229_));
 sky130_fd_sc_hd__xnor2_2 _28883_ (.A(_00228_),
    .B(_00229_),
    .Y(_00231_));
 sky130_fd_sc_hd__nor2_2 _28884_ (.A(_14988_),
    .B(_15173_),
    .Y(_00232_));
 sky130_fd_sc_hd__xnor2_2 _28885_ (.A(_00231_),
    .B(_00232_),
    .Y(_00233_));
 sky130_fd_sc_hd__or3_2 _28886_ (.A(_14612_),
    .B(_17696_),
    .C(_18792_),
    .X(_00234_));
 sky130_fd_sc_hd__o21ai_2 _28887_ (.A1(_14612_),
    .A2(_17696_),
    .B1(_18792_),
    .Y(_00235_));
 sky130_fd_sc_hd__nand2_2 _28888_ (.A(_00234_),
    .B(_00235_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_2 _28889_ (.A(_14392_),
    .B(_17460_),
    .Y(_00237_));
 sky130_fd_sc_hd__xnor2_2 _28890_ (.A(_00236_),
    .B(_00237_),
    .Y(_00238_));
 sky130_fd_sc_hd__or3_2 _28891_ (.A(_18791_),
    .B(_18180_),
    .C(_18792_),
    .X(_00239_));
 sky130_fd_sc_hd__o21a_2 _28892_ (.A1(_18794_),
    .A2(_18795_),
    .B1(_00239_),
    .X(_00240_));
 sky130_fd_sc_hd__xnor2_2 _28893_ (.A(_00238_),
    .B(_00240_),
    .Y(_00242_));
 sky130_fd_sc_hd__xor2_2 _28894_ (.A(_00233_),
    .B(_00242_),
    .X(_00243_));
 sky130_fd_sc_hd__o21ai_2 _28895_ (.A1(_00226_),
    .A2(_00227_),
    .B1(_00243_),
    .Y(_00244_));
 sky130_fd_sc_hd__or3_2 _28896_ (.A(_00226_),
    .B(_00227_),
    .C(_00243_),
    .X(_00245_));
 sky130_fd_sc_hd__and2_2 _28897_ (.A(_00244_),
    .B(_00245_),
    .X(_00246_));
 sky130_fd_sc_hd__xnor2_2 _28898_ (.A(_00225_),
    .B(_00246_),
    .Y(_00247_));
 sky130_fd_sc_hd__a21bo_2 _28899_ (.A1(_18805_),
    .A2(_18807_),
    .B1_N(_18804_),
    .X(_00248_));
 sky130_fd_sc_hd__a31o_2 _28900_ (.A1(_15887_),
    .A2(_17702_),
    .A3(_18814_),
    .B1(_18813_),
    .X(_00249_));
 sky130_fd_sc_hd__nor2_2 _28901_ (.A(_12850_),
    .B(_16999_),
    .Y(_00250_));
 sky130_fd_sc_hd__or3b_2 _28902_ (.A(_12848_),
    .B(_17007_),
    .C_N(_00250_),
    .X(_00251_));
 sky130_fd_sc_hd__a22o_2 _28903_ (.A1(_12846_),
    .A2(_16680_),
    .B1(_17003_),
    .B2(_14636_),
    .X(_00253_));
 sky130_fd_sc_hd__nand2_2 _28904_ (.A(_00251_),
    .B(_00253_),
    .Y(_00254_));
 sky130_fd_sc_hd__buf_1 _28905_ (.A(_16988_),
    .X(_00255_));
 sky130_fd_sc_hd__nor2_2 _28906_ (.A(_14625_),
    .B(_00255_),
    .Y(_00256_));
 sky130_fd_sc_hd__xnor2_2 _28907_ (.A(_00254_),
    .B(_00256_),
    .Y(_00257_));
 sky130_fd_sc_hd__xor2_2 _28908_ (.A(_00249_),
    .B(_00257_),
    .X(_00258_));
 sky130_fd_sc_hd__and2_2 _28909_ (.A(_00248_),
    .B(_00258_),
    .X(_00259_));
 sky130_fd_sc_hd__nor2_2 _28910_ (.A(_00248_),
    .B(_00258_),
    .Y(_00260_));
 sky130_fd_sc_hd__nor2_2 _28911_ (.A(_00259_),
    .B(_00260_),
    .Y(_00261_));
 sky130_fd_sc_hd__nand2_2 _28912_ (.A(_15887_),
    .B(_18209_),
    .Y(_00262_));
 sky130_fd_sc_hd__and4_2 _28913_ (.A(_14649_),
    .B(_12243_),
    .C(_18205_),
    .D(_18203_),
    .X(_00264_));
 sky130_fd_sc_hd__o22a_2 _28914_ (.A1(_14978_),
    .A2(_18443_),
    .B1(_18211_),
    .B2(_15650_),
    .X(_00265_));
 sky130_fd_sc_hd__nor2_2 _28915_ (.A(_00264_),
    .B(_00265_),
    .Y(_00266_));
 sky130_fd_sc_hd__xnor2_2 _28916_ (.A(_00262_),
    .B(_00266_),
    .Y(_00267_));
 sky130_fd_sc_hd__nor2_2 _28917_ (.A(_18822_),
    .B(_18823_),
    .Y(_00268_));
 sky130_fd_sc_hd__and3_2 _28918_ (.A(_11381_),
    .B(_18457_),
    .C(_00268_),
    .X(_00269_));
 sky130_fd_sc_hd__nor3_2 _28919_ (.A(_11793_),
    .B(_18211_),
    .C(_18825_),
    .Y(_00270_));
 sky130_fd_sc_hd__buf_1 _28920_ (.A(_18456_),
    .X(_00271_));
 sky130_fd_sc_hd__nor2_2 _28921_ (.A(_11793_),
    .B(_00271_),
    .Y(_00272_));
 sky130_fd_sc_hd__or3_2 _28922_ (.A(_11575_),
    .B(_18822_),
    .C(_18823_),
    .X(_00273_));
 sky130_fd_sc_hd__nand2_2 _28923_ (.A(iX[26]),
    .B(iX[58]),
    .Y(_00275_));
 sky130_fd_sc_hd__or2_2 _28924_ (.A(iX[26]),
    .B(iX[58]),
    .X(_00276_));
 sky130_fd_sc_hd__nand2_2 _28925_ (.A(_00275_),
    .B(_00276_),
    .Y(_00277_));
 sky130_fd_sc_hd__a311oi_2 _28926_ (.A1(_18451_),
    .A2(_18454_),
    .A3(_18819_),
    .B1(_00277_),
    .C1(_18818_),
    .Y(_00278_));
 sky130_fd_sc_hd__a21o_2 _28927_ (.A1(_18451_),
    .A2(_18819_),
    .B1(_18818_),
    .X(_00279_));
 sky130_fd_sc_hd__o211a_2 _28928_ (.A1(_18454_),
    .A2(_18818_),
    .B1(_00277_),
    .C1(_00279_),
    .X(_00280_));
 sky130_fd_sc_hd__or3_2 _28929_ (.A(_11565_),
    .B(_00278_),
    .C(_00280_),
    .X(_00281_));
 sky130_fd_sc_hd__xor2_2 _28930_ (.A(_00273_),
    .B(_00281_),
    .X(_00282_));
 sky130_fd_sc_hd__xnor2_2 _28931_ (.A(_00272_),
    .B(_00282_),
    .Y(_00283_));
 sky130_fd_sc_hd__o21bai_2 _28932_ (.A1(_00269_),
    .A2(_00270_),
    .B1_N(_00283_),
    .Y(_00284_));
 sky130_fd_sc_hd__or3b_2 _28933_ (.A(_00269_),
    .B(_00270_),
    .C_N(_00283_),
    .X(_00286_));
 sky130_fd_sc_hd__and3_2 _28934_ (.A(_00267_),
    .B(_00284_),
    .C(_00286_),
    .X(_00287_));
 sky130_fd_sc_hd__a21oi_2 _28935_ (.A1(_00284_),
    .A2(_00286_),
    .B1(_00267_),
    .Y(_00288_));
 sky130_fd_sc_hd__or2_4 _28936_ (.A(_00287_),
    .B(_00288_),
    .X(_00289_));
 sky130_fd_sc_hd__and2_2 _28937_ (.A(_18826_),
    .B(_18827_),
    .X(_00290_));
 sky130_fd_sc_hd__a21oi_2 _28938_ (.A1(_18816_),
    .A2(_18828_),
    .B1(_00290_),
    .Y(_00291_));
 sky130_fd_sc_hd__xor2_2 _28939_ (.A(_00289_),
    .B(_00291_),
    .X(_00292_));
 sky130_fd_sc_hd__xnor2_2 _28940_ (.A(_00261_),
    .B(_00292_),
    .Y(_00293_));
 sky130_fd_sc_hd__and2b_2 _28941_ (.A_N(_18829_),
    .B(_18830_),
    .X(_00294_));
 sky130_fd_sc_hd__and2b_2 _28942_ (.A_N(_18811_),
    .B(_18832_),
    .X(_00295_));
 sky130_fd_sc_hd__nor2_2 _28943_ (.A(_00294_),
    .B(_00295_),
    .Y(_00297_));
 sky130_fd_sc_hd__xor2_2 _28944_ (.A(_00293_),
    .B(_00297_),
    .X(_00298_));
 sky130_fd_sc_hd__xor2_2 _28945_ (.A(_00247_),
    .B(_00298_),
    .X(_00299_));
 sky130_fd_sc_hd__and2b_2 _28946_ (.A_N(_18801_),
    .B(_18835_),
    .X(_00300_));
 sky130_fd_sc_hd__a21oi_2 _28947_ (.A1(_18833_),
    .A2(_18834_),
    .B1(_00300_),
    .Y(_00301_));
 sky130_fd_sc_hd__xnor2_2 _28948_ (.A(_00299_),
    .B(_00301_),
    .Y(_00302_));
 sky130_fd_sc_hd__xnor2_2 _28949_ (.A(_00223_),
    .B(_00302_),
    .Y(_00303_));
 sky130_fd_sc_hd__and2b_2 _28950_ (.A_N(_18837_),
    .B(_18836_),
    .X(_00304_));
 sky130_fd_sc_hd__a21o_2 _28951_ (.A1(_18780_),
    .A2(_18838_),
    .B1(_00304_),
    .X(_00305_));
 sky130_fd_sc_hd__xor2_2 _28952_ (.A(_00303_),
    .B(_00305_),
    .X(_00306_));
 sky130_fd_sc_hd__xnor2_2 _28953_ (.A(_00178_),
    .B(_00306_),
    .Y(_00308_));
 sky130_fd_sc_hd__or2b_2 _28954_ (.A(_18839_),
    .B_N(_18840_),
    .X(_00309_));
 sky130_fd_sc_hd__o21ai_2 _28955_ (.A1(_18745_),
    .A2(_18841_),
    .B1(_00309_),
    .Y(_00310_));
 sky130_fd_sc_hd__xnor2_2 _28956_ (.A(_00308_),
    .B(_00310_),
    .Y(_00311_));
 sky130_fd_sc_hd__xor2_2 _28957_ (.A(_00146_),
    .B(_00311_),
    .X(_00312_));
 sky130_fd_sc_hd__xnor2_2 _28958_ (.A(_00144_),
    .B(_00312_),
    .Y(_00313_));
 sky130_fd_sc_hd__xnor2_2 _28959_ (.A(_00140_),
    .B(_00313_),
    .Y(_00314_));
 sky130_fd_sc_hd__nor2_2 _28960_ (.A(_18497_),
    .B(_18850_),
    .Y(_00315_));
 sky130_fd_sc_hd__a21o_2 _28961_ (.A1(_18716_),
    .A2(_00315_),
    .B1(_18849_),
    .X(_00316_));
 sky130_fd_sc_hd__xnor2_2 _28962_ (.A(_00314_),
    .B(_00316_),
    .Y(_00317_));
 sky130_fd_sc_hd__nand2_2 _28963_ (.A(_18922_),
    .B(_18923_),
    .Y(_00319_));
 sky130_fd_sc_hd__or3_2 _28964_ (.A(_18924_),
    .B(_00031_),
    .C(_00032_),
    .X(_00320_));
 sky130_fd_sc_hd__nor2_2 _28965_ (.A(_18894_),
    .B(_18921_),
    .Y(_00321_));
 sky130_fd_sc_hd__or2b_2 _28966_ (.A(_18867_),
    .B_N(_18866_),
    .X(_00322_));
 sky130_fd_sc_hd__and4_2 _28967_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[55]),
    .D(iX[56]),
    .X(_00323_));
 sky130_fd_sc_hd__a22oi_2 _28968_ (.A1(iY[35]),
    .A2(iX[55]),
    .B1(iX[56]),
    .B2(iY[34]),
    .Y(_00324_));
 sky130_fd_sc_hd__nor2_2 _28969_ (.A(_00323_),
    .B(_00324_),
    .Y(_00325_));
 sky130_fd_sc_hd__nand2_2 _28970_ (.A(iY[33]),
    .B(iX[57]),
    .Y(_00326_));
 sky130_fd_sc_hd__xnor2_2 _28971_ (.A(_00325_),
    .B(_00326_),
    .Y(_00327_));
 sky130_fd_sc_hd__o21ba_2 _28972_ (.A1(_18862_),
    .A2(_18865_),
    .B1_N(_18861_),
    .X(_00328_));
 sky130_fd_sc_hd__xnor2_2 _28973_ (.A(_00327_),
    .B(_00328_),
    .Y(_00330_));
 sky130_fd_sc_hd__and4_2 _28974_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[54]),
    .D(iX[58]),
    .X(_00331_));
 sky130_fd_sc_hd__a22oi_2 _28975_ (.A1(iY[36]),
    .A2(iX[54]),
    .B1(iX[58]),
    .B2(iY[32]),
    .Y(_00332_));
 sky130_fd_sc_hd__nor2_2 _28976_ (.A(_00331_),
    .B(_00332_),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_2 _28977_ (.A(iY[37]),
    .B(iX[53]),
    .Y(_00334_));
 sky130_fd_sc_hd__xnor2_2 _28978_ (.A(_00333_),
    .B(_00334_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_2 _28979_ (.A(_00330_),
    .B(_00335_),
    .Y(_00336_));
 sky130_fd_sc_hd__or2_2 _28980_ (.A(_00330_),
    .B(_00335_),
    .X(_00337_));
 sky130_fd_sc_hd__nand2_2 _28981_ (.A(_00336_),
    .B(_00337_),
    .Y(_00338_));
 sky130_fd_sc_hd__a21o_2 _28982_ (.A1(_00322_),
    .A2(_18874_),
    .B1(_00338_),
    .X(_00339_));
 sky130_fd_sc_hd__nand3_2 _28983_ (.A(_00322_),
    .B(_18874_),
    .C(_00338_),
    .Y(_00341_));
 sky130_fd_sc_hd__o21ba_2 _28984_ (.A1(_18883_),
    .A2(_18885_),
    .B1_N(_18882_),
    .X(_00342_));
 sky130_fd_sc_hd__o21ba_2 _28985_ (.A1(_18870_),
    .A2(_18872_),
    .B1_N(_18869_),
    .X(_00343_));
 sky130_fd_sc_hd__and4_2 _28986_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[51]),
    .D(iX[52]),
    .X(_00344_));
 sky130_fd_sc_hd__a22oi_2 _28987_ (.A1(iY[39]),
    .A2(iX[51]),
    .B1(iX[52]),
    .B2(iY[38]),
    .Y(_00345_));
 sky130_fd_sc_hd__nor2_2 _28988_ (.A(_00344_),
    .B(_00345_),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_2 _28989_ (.A(iY[40]),
    .B(iX[50]),
    .Y(_00347_));
 sky130_fd_sc_hd__xnor2_2 _28990_ (.A(_00346_),
    .B(_00347_),
    .Y(_00348_));
 sky130_fd_sc_hd__xnor2_2 _28991_ (.A(_00343_),
    .B(_00348_),
    .Y(_00349_));
 sky130_fd_sc_hd__xnor2_2 _28992_ (.A(_00342_),
    .B(_00349_),
    .Y(_00350_));
 sky130_fd_sc_hd__and3_2 _28993_ (.A(_00339_),
    .B(_00341_),
    .C(_00350_),
    .X(_00352_));
 sky130_fd_sc_hd__a21oi_2 _28994_ (.A1(_00339_),
    .A2(_00341_),
    .B1(_00350_),
    .Y(_00353_));
 sky130_fd_sc_hd__nor2_2 _28995_ (.A(_00352_),
    .B(_00353_),
    .Y(_00354_));
 sky130_fd_sc_hd__nand2_2 _28996_ (.A(_18878_),
    .B(_18890_),
    .Y(_00355_));
 sky130_fd_sc_hd__xnor2_2 _28997_ (.A(_00354_),
    .B(_00355_),
    .Y(_00356_));
 sky130_fd_sc_hd__and2b_2 _28998_ (.A_N(_18911_),
    .B(_18910_),
    .X(_00357_));
 sky130_fd_sc_hd__or2b_2 _28999_ (.A(_18881_),
    .B_N(_18887_),
    .X(_00358_));
 sky130_fd_sc_hd__or2b_2 _29000_ (.A(_18880_),
    .B_N(_18888_),
    .X(_00359_));
 sky130_fd_sc_hd__and4_2 _29001_ (.A(iY[44]),
    .B(iX[45]),
    .C(iY[45]),
    .D(iX[46]),
    .X(_00360_));
 sky130_fd_sc_hd__a22oi_2 _29002_ (.A1(iX[45]),
    .A2(iY[45]),
    .B1(iX[46]),
    .B2(iY[44]),
    .Y(_00361_));
 sky130_fd_sc_hd__nor2_2 _29003_ (.A(_00360_),
    .B(_00361_),
    .Y(_00363_));
 sky130_fd_sc_hd__nand2_2 _29004_ (.A(iX[44]),
    .B(iY[46]),
    .Y(_00364_));
 sky130_fd_sc_hd__xnor2_2 _29005_ (.A(_00363_),
    .B(_00364_),
    .Y(_00365_));
 sky130_fd_sc_hd__and4_2 _29006_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[48]),
    .D(iX[49]),
    .X(_00366_));
 sky130_fd_sc_hd__a22oi_2 _29007_ (.A1(iY[42]),
    .A2(iX[48]),
    .B1(iX[49]),
    .B2(iY[41]),
    .Y(_00367_));
 sky130_fd_sc_hd__nor2_2 _29008_ (.A(_00366_),
    .B(_00367_),
    .Y(_00368_));
 sky130_fd_sc_hd__nand2_2 _29009_ (.A(iY[43]),
    .B(iX[47]),
    .Y(_00369_));
 sky130_fd_sc_hd__xnor2_2 _29010_ (.A(_00368_),
    .B(_00369_),
    .Y(_00370_));
 sky130_fd_sc_hd__o21ai_2 _29011_ (.A1(_18905_),
    .A2(_18907_),
    .B1(_00370_),
    .Y(_00371_));
 sky130_fd_sc_hd__or3_2 _29012_ (.A(_18905_),
    .B(_18907_),
    .C(_00370_),
    .X(_00372_));
 sky130_fd_sc_hd__and2_2 _29013_ (.A(_00371_),
    .B(_00372_),
    .X(_00374_));
 sky130_fd_sc_hd__xnor2_2 _29014_ (.A(_00365_),
    .B(_00374_),
    .Y(_00375_));
 sky130_fd_sc_hd__a21oi_2 _29015_ (.A1(_00358_),
    .A2(_00359_),
    .B1(_00375_),
    .Y(_00376_));
 sky130_fd_sc_hd__inv_2 _29016_ (.A(_00376_),
    .Y(_00377_));
 sky130_fd_sc_hd__nand3_2 _29017_ (.A(_00358_),
    .B(_00359_),
    .C(_00375_),
    .Y(_00378_));
 sky130_fd_sc_hd__o211a_2 _29018_ (.A1(_00357_),
    .A2(_18913_),
    .B1(_00377_),
    .C1(_00378_),
    .X(_00379_));
 sky130_fd_sc_hd__a211o_2 _29019_ (.A1(_00377_),
    .A2(_00378_),
    .B1(_00357_),
    .C1(_18913_),
    .X(_00380_));
 sky130_fd_sc_hd__or3b_2 _29020_ (.A(_00356_),
    .B(_00379_),
    .C_N(_00380_),
    .X(_00381_));
 sky130_fd_sc_hd__inv_2 _29021_ (.A(_00379_),
    .Y(_00382_));
 sky130_fd_sc_hd__a21bo_2 _29022_ (.A1(_00382_),
    .A2(_00380_),
    .B1_N(_00356_),
    .X(_00383_));
 sky130_fd_sc_hd__o211a_2 _29023_ (.A1(_18892_),
    .A2(_00321_),
    .B1(_00381_),
    .C1(_00383_),
    .X(_00385_));
 sky130_fd_sc_hd__a211oi_2 _29024_ (.A1(_00381_),
    .A2(_00383_),
    .B1(_18892_),
    .C1(_00321_),
    .Y(_00386_));
 sky130_fd_sc_hd__a21o_2 _29025_ (.A1(_00012_),
    .A2(_18604_),
    .B1(_00023_),
    .X(_00387_));
 sky130_fd_sc_hd__and4_2 _29026_ (.A(iX[36]),
    .B(iX[37]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_00388_));
 sky130_fd_sc_hd__a22oi_2 _29027_ (.A1(iX[37]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[36]),
    .Y(_00389_));
 sky130_fd_sc_hd__nor2_2 _29028_ (.A(_00388_),
    .B(_00389_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_2 _29029_ (.A(iX[35]),
    .B(iY[55]),
    .Y(_00391_));
 sky130_fd_sc_hd__xnor2_2 _29030_ (.A(_00390_),
    .B(_00391_),
    .Y(_00392_));
 sky130_fd_sc_hd__and4_2 _29031_ (.A(iX[39]),
    .B(iX[40]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_00393_));
 sky130_fd_sc_hd__a22oi_2 _29032_ (.A1(iX[40]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[39]),
    .Y(_00394_));
 sky130_fd_sc_hd__nor2_2 _29033_ (.A(_00393_),
    .B(_00394_),
    .Y(_00396_));
 sky130_fd_sc_hd__nand2_2 _29034_ (.A(iX[38]),
    .B(iY[52]),
    .Y(_00397_));
 sky130_fd_sc_hd__xnor2_2 _29035_ (.A(_00396_),
    .B(_00397_),
    .Y(_00398_));
 sky130_fd_sc_hd__o21ba_2 _29036_ (.A1(_00002_),
    .A2(_00004_),
    .B1_N(_00001_),
    .X(_00399_));
 sky130_fd_sc_hd__xnor2_2 _29037_ (.A(_00398_),
    .B(_00399_),
    .Y(_00400_));
 sky130_fd_sc_hd__and2_2 _29038_ (.A(_00392_),
    .B(_00400_),
    .X(_00401_));
 sky130_fd_sc_hd__nor2_2 _29039_ (.A(_00392_),
    .B(_00400_),
    .Y(_00402_));
 sky130_fd_sc_hd__or2_2 _29040_ (.A(_00401_),
    .B(_00402_),
    .X(_00403_));
 sky130_fd_sc_hd__or3_2 _29041_ (.A(_00013_),
    .B(_00016_),
    .C(_00017_),
    .X(_00404_));
 sky130_fd_sc_hd__o21ba_2 _29042_ (.A1(_18901_),
    .A2(_18903_),
    .B1_N(_18900_),
    .X(_00405_));
 sky130_fd_sc_hd__and4_2 _29043_ (.A(iX[42]),
    .B(iX[43]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_00407_));
 sky130_fd_sc_hd__a22oi_2 _29044_ (.A1(iX[43]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[42]),
    .Y(_00408_));
 sky130_fd_sc_hd__and4bb_2 _29045_ (.A_N(_00407_),
    .B_N(_00408_),
    .C(iX[41]),
    .D(iY[49]),
    .X(_00409_));
 sky130_fd_sc_hd__o2bb2a_2 _29046_ (.A1_N(iX[41]),
    .A2_N(iY[49]),
    .B1(_00407_),
    .B2(_00408_),
    .X(_00410_));
 sky130_fd_sc_hd__nor2_2 _29047_ (.A(_00409_),
    .B(_00410_),
    .Y(_00411_));
 sky130_fd_sc_hd__xnor2_2 _29048_ (.A(_00405_),
    .B(_00411_),
    .Y(_00412_));
 sky130_fd_sc_hd__o21ai_2 _29049_ (.A1(_00014_),
    .A2(_00016_),
    .B1(_00412_),
    .Y(_00413_));
 sky130_fd_sc_hd__or3_2 _29050_ (.A(_00014_),
    .B(_00016_),
    .C(_00412_),
    .X(_00414_));
 sky130_fd_sc_hd__nand2_2 _29051_ (.A(_00413_),
    .B(_00414_),
    .Y(_00415_));
 sky130_fd_sc_hd__a21oi_2 _29052_ (.A1(_00404_),
    .A2(_00020_),
    .B1(_00415_),
    .Y(_00416_));
 sky130_fd_sc_hd__and3_2 _29053_ (.A(_00404_),
    .B(_00020_),
    .C(_00415_),
    .X(_00418_));
 sky130_fd_sc_hd__nor3_2 _29054_ (.A(_00403_),
    .B(_00416_),
    .C(_00418_),
    .Y(_00419_));
 sky130_fd_sc_hd__o21a_2 _29055_ (.A1(_00416_),
    .A2(_00418_),
    .B1(_00403_),
    .X(_00420_));
 sky130_fd_sc_hd__a211oi_2 _29056_ (.A1(_18916_),
    .A2(_18918_),
    .B1(_00419_),
    .C1(_00420_),
    .Y(_00421_));
 sky130_fd_sc_hd__o211a_2 _29057_ (.A1(_00419_),
    .A2(_00420_),
    .B1(_18916_),
    .C1(_18918_),
    .X(_00422_));
 sky130_fd_sc_hd__a211oi_2 _29058_ (.A1(_00387_),
    .A2(_00026_),
    .B1(_00421_),
    .C1(_00422_),
    .Y(_00423_));
 sky130_fd_sc_hd__o211a_2 _29059_ (.A1(_00421_),
    .A2(_00422_),
    .B1(_00387_),
    .C1(_00026_),
    .X(_00424_));
 sky130_fd_sc_hd__nor4_2 _29060_ (.A(_00385_),
    .B(_00386_),
    .C(_00423_),
    .D(_00424_),
    .Y(_00425_));
 sky130_fd_sc_hd__o22a_2 _29061_ (.A1(_00385_),
    .A2(_00386_),
    .B1(_00423_),
    .B2(_00424_),
    .X(_00426_));
 sky130_fd_sc_hd__a211oi_2 _29062_ (.A1(_00319_),
    .A2(_00320_),
    .B1(_00425_),
    .C1(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__o211a_2 _29063_ (.A1(_00425_),
    .A2(_00426_),
    .B1(_00319_),
    .C1(_00320_),
    .X(_00429_));
 sky130_fd_sc_hd__or2_2 _29064_ (.A(_00028_),
    .B(_00031_),
    .X(_00430_));
 sky130_fd_sc_hd__or2b_2 _29065_ (.A(_00006_),
    .B_N(_00005_),
    .X(_00431_));
 sky130_fd_sc_hd__o21ba_2 _29066_ (.A1(_18926_),
    .A2(_18928_),
    .B1_N(_18925_),
    .X(_00432_));
 sky130_fd_sc_hd__and4_2 _29067_ (.A(iX[33]),
    .B(iX[34]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_00433_));
 sky130_fd_sc_hd__a22oi_2 _29068_ (.A1(iX[34]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[33]),
    .Y(_00434_));
 sky130_fd_sc_hd__nor2_2 _29069_ (.A(_00433_),
    .B(_00434_),
    .Y(_00435_));
 sky130_fd_sc_hd__nand2_2 _29070_ (.A(iX[32]),
    .B(iY[58]),
    .Y(_00436_));
 sky130_fd_sc_hd__xnor2_2 _29071_ (.A(_00435_),
    .B(_00436_),
    .Y(_00437_));
 sky130_fd_sc_hd__xnor2_2 _29072_ (.A(_00432_),
    .B(_00437_),
    .Y(_00438_));
 sky130_fd_sc_hd__xnor2_2 _29073_ (.A(_00042_),
    .B(_00438_),
    .Y(_00440_));
 sky130_fd_sc_hd__a21oi_2 _29074_ (.A1(_00431_),
    .A2(_00008_),
    .B1(_00440_),
    .Y(_00441_));
 sky130_fd_sc_hd__and3_2 _29075_ (.A(_00431_),
    .B(_00008_),
    .C(_00440_),
    .X(_00442_));
 sky130_fd_sc_hd__nor2_2 _29076_ (.A(_00441_),
    .B(_00442_),
    .Y(_00443_));
 sky130_fd_sc_hd__xnor2_2 _29077_ (.A(_00045_),
    .B(_00443_),
    .Y(_00444_));
 sky130_fd_sc_hd__a21o_2 _29078_ (.A1(_00048_),
    .A2(_00051_),
    .B1(_00444_),
    .X(_00445_));
 sky130_fd_sc_hd__nand3_2 _29079_ (.A(_00048_),
    .B(_00051_),
    .C(_00444_),
    .Y(_00446_));
 sky130_fd_sc_hd__nand2_2 _29080_ (.A(_00445_),
    .B(_00446_),
    .Y(_00447_));
 sky130_fd_sc_hd__xnor2_2 _29081_ (.A(_00430_),
    .B(_00447_),
    .Y(_00448_));
 sky130_fd_sc_hd__nor2_2 _29082_ (.A(_00054_),
    .B(_00448_),
    .Y(_00449_));
 sky130_fd_sc_hd__and2_2 _29083_ (.A(_00054_),
    .B(_00448_),
    .X(_00451_));
 sky130_fd_sc_hd__or2_2 _29084_ (.A(_00449_),
    .B(_00451_),
    .X(_00452_));
 sky130_fd_sc_hd__or3_2 _29085_ (.A(_00427_),
    .B(_00429_),
    .C(_00452_),
    .X(_00453_));
 sky130_fd_sc_hd__o21ai_2 _29086_ (.A1(_00427_),
    .A2(_00429_),
    .B1(_00452_),
    .Y(_00454_));
 sky130_fd_sc_hd__o211ai_2 _29087_ (.A1(_00036_),
    .A2(_00062_),
    .B1(_00453_),
    .C1(_00454_),
    .Y(_00455_));
 sky130_fd_sc_hd__a211o_2 _29088_ (.A1(_00453_),
    .A2(_00454_),
    .B1(_00036_),
    .C1(_00062_),
    .X(_00456_));
 sky130_fd_sc_hd__nand2_2 _29089_ (.A(_00455_),
    .B(_00456_),
    .Y(_00457_));
 sky130_fd_sc_hd__a21oi_2 _29090_ (.A1(_00038_),
    .A2(_00060_),
    .B1(_00058_),
    .Y(_00458_));
 sky130_fd_sc_hd__xnor2_2 _29091_ (.A(_00457_),
    .B(_00458_),
    .Y(_00459_));
 sky130_fd_sc_hd__a21oi_2 _29092_ (.A1(_00065_),
    .A2(_00068_),
    .B1(_00459_),
    .Y(_00460_));
 sky130_fd_sc_hd__and3_2 _29093_ (.A(_00065_),
    .B(_00068_),
    .C(_00459_),
    .X(_00462_));
 sky130_fd_sc_hd__nor2_2 _29094_ (.A(_00460_),
    .B(_00462_),
    .Y(_00463_));
 sky130_fd_sc_hd__xnor2_2 _29095_ (.A(_00070_),
    .B(_00463_),
    .Y(_00464_));
 sky130_fd_sc_hd__nand2_2 _29096_ (.A(_18645_),
    .B(_00074_),
    .Y(_00465_));
 sky130_fd_sc_hd__a31o_2 _29097_ (.A1(_18502_),
    .A2(_18504_),
    .A3(_18507_),
    .B1(_00465_),
    .X(_00466_));
 sky130_fd_sc_hd__a21oi_2 _29098_ (.A1(_18643_),
    .A2(_00074_),
    .B1(_00072_),
    .Y(_00467_));
 sky130_fd_sc_hd__and2_2 _29099_ (.A(_00466_),
    .B(_00467_),
    .X(_00468_));
 sky130_fd_sc_hd__xnor2_2 _29100_ (.A(_00464_),
    .B(_00468_),
    .Y(_00469_));
 sky130_fd_sc_hd__xor2_2 _29101_ (.A(_00317_),
    .B(_00469_),
    .X(_00470_));
 sky130_fd_sc_hd__xnor2_2 _29102_ (.A(_10382_),
    .B(_00470_),
    .Y(_00471_));
 sky130_fd_sc_hd__a21oi_2 _29103_ (.A1(_00139_),
    .A2(_00080_),
    .B1(_00471_),
    .Y(_00473_));
 sky130_fd_sc_hd__nand3_2 _29104_ (.A(_00139_),
    .B(_00080_),
    .C(_00471_),
    .Y(_00474_));
 sky130_fd_sc_hd__or2b_2 _29105_ (.A(_00473_),
    .B_N(_00474_),
    .X(_00475_));
 sky130_fd_sc_hd__or3_4 _29106_ (.A(_18652_),
    .B(_00084_),
    .C(_00085_),
    .X(_00476_));
 sky130_fd_sc_hd__a2111o_2 _29107_ (.A1(_17877_),
    .A2(_18654_),
    .B1(_00476_),
    .C1(_18259_),
    .D1(_18655_),
    .X(_00477_));
 sky130_fd_sc_hd__inv_2 _29108_ (.A(_00087_),
    .Y(_00478_));
 sky130_fd_sc_hd__o21bai_2 _29109_ (.A1(_00478_),
    .A2(_00084_),
    .B1_N(_00085_),
    .Y(_00479_));
 sky130_fd_sc_hd__nand2_2 _29110_ (.A(_00477_),
    .B(_00479_),
    .Y(_00480_));
 sky130_fd_sc_hd__xnor2_2 _29111_ (.A(_00475_),
    .B(_00480_),
    .Y(_00481_));
 sky130_fd_sc_hd__and2_2 _29112_ (.A(_00138_),
    .B(_00481_),
    .X(_00482_));
 sky130_fd_sc_hd__nor2_2 _29113_ (.A(_00138_),
    .B(_00481_),
    .Y(_00484_));
 sky130_fd_sc_hd__nor2_2 _29114_ (.A(_00482_),
    .B(_00484_),
    .Y(_00485_));
 sky130_fd_sc_hd__o21a_2 _29115_ (.A1(_00097_),
    .A2(_00100_),
    .B1(_00485_),
    .X(_00486_));
 sky130_fd_sc_hd__nor3_2 _29116_ (.A(_00485_),
    .B(_00097_),
    .C(_00100_),
    .Y(_00487_));
 sky130_fd_sc_hd__nor2_2 _29117_ (.A(_00486_),
    .B(_00487_),
    .Y(oO[58]));
 sky130_fd_sc_hd__and3_2 _29118_ (.A(_18302_),
    .B(_18698_),
    .C(_00125_),
    .X(_00488_));
 sky130_fd_sc_hd__and3_2 _29119_ (.A(_18694_),
    .B(_18695_),
    .C(_00125_),
    .X(_00489_));
 sky130_fd_sc_hd__nor2_2 _29120_ (.A(_00106_),
    .B(_00107_),
    .Y(_00490_));
 sky130_fd_sc_hd__nand2_2 _29121_ (.A(iY[29]),
    .B(iX[31]),
    .Y(_00491_));
 sky130_fd_sc_hd__a22o_2 _29122_ (.A1(iY[29]),
    .A2(iX[30]),
    .B1(iX[31]),
    .B2(iY[28]),
    .X(_00492_));
 sky130_fd_sc_hd__o21a_2 _29123_ (.A1(_00103_),
    .A2(_00491_),
    .B1(_00492_),
    .X(_00494_));
 sky130_fd_sc_hd__o21a_2 _29124_ (.A1(_00105_),
    .A2(_00490_),
    .B1(_00494_),
    .X(_00495_));
 sky130_fd_sc_hd__nor3_2 _29125_ (.A(_00105_),
    .B(_00490_),
    .C(_00494_),
    .Y(_00496_));
 sky130_fd_sc_hd__nor2_2 _29126_ (.A(_00495_),
    .B(_00496_),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_2 _29127_ (.A(iX[29]),
    .B(iY[30]),
    .Y(_00498_));
 sky130_fd_sc_hd__xor2_2 _29128_ (.A(_00497_),
    .B(_00498_),
    .X(_00499_));
 sky130_fd_sc_hd__and2b_2 _29129_ (.A_N(_00110_),
    .B(_00108_),
    .X(_00500_));
 sky130_fd_sc_hd__a31oi_2 _29130_ (.A1(iX[28]),
    .A2(iY[30]),
    .A3(_00111_),
    .B1(_00500_),
    .Y(_00501_));
 sky130_fd_sc_hd__xnor2_2 _29131_ (.A(_00499_),
    .B(_00501_),
    .Y(_00502_));
 sky130_fd_sc_hd__nand2_2 _29132_ (.A(iX[28]),
    .B(iY[31]),
    .Y(_00503_));
 sky130_fd_sc_hd__and2_2 _29133_ (.A(_00502_),
    .B(_00503_),
    .X(_00505_));
 sky130_fd_sc_hd__nor2_2 _29134_ (.A(_00502_),
    .B(_00503_),
    .Y(_00506_));
 sky130_fd_sc_hd__nor2_2 _29135_ (.A(_00505_),
    .B(_00506_),
    .Y(_00507_));
 sky130_fd_sc_hd__a21oi_2 _29136_ (.A1(_00123_),
    .A2(_00124_),
    .B1(_00507_),
    .Y(_00508_));
 sky130_fd_sc_hd__and3_2 _29137_ (.A(_00123_),
    .B(_00124_),
    .C(_00507_),
    .X(_00509_));
 sky130_fd_sc_hd__and3_2 _29138_ (.A(_00118_),
    .B(_00119_),
    .C(_00507_),
    .X(_00510_));
 sky130_fd_sc_hd__a211oi_2 _29139_ (.A1(_00121_),
    .A2(_00508_),
    .B1(_00509_),
    .C1(_00510_),
    .Y(_00511_));
 sky130_fd_sc_hd__nand2_2 _29140_ (.A(_00489_),
    .B(_00511_),
    .Y(_00512_));
 sky130_fd_sc_hd__or2_2 _29141_ (.A(_00489_),
    .B(_00511_),
    .X(_00513_));
 sky130_fd_sc_hd__nand2_2 _29142_ (.A(_00512_),
    .B(_00513_),
    .Y(_00514_));
 sky130_fd_sc_hd__a31o_2 _29143_ (.A1(iX[27]),
    .A2(iY[31]),
    .A3(_00116_),
    .B1(_00114_),
    .X(_00516_));
 sky130_fd_sc_hd__xnor2_2 _29144_ (.A(_00514_),
    .B(_00516_),
    .Y(_00517_));
 sky130_fd_sc_hd__o21a_2 _29145_ (.A1(_00128_),
    .A2(_00488_),
    .B1(_00517_),
    .X(_00518_));
 sky130_fd_sc_hd__nor3_2 _29146_ (.A(_00128_),
    .B(_00517_),
    .C(_00488_),
    .Y(_00519_));
 sky130_fd_sc_hd__or2_2 _29147_ (.A(_00518_),
    .B(_00519_),
    .X(_00520_));
 sky130_fd_sc_hd__nor2_2 _29148_ (.A(_00133_),
    .B(_00136_),
    .Y(_00521_));
 sky130_fd_sc_hd__xnor2_2 _29149_ (.A(_00520_),
    .B(_00521_),
    .Y(_00522_));
 sky130_fd_sc_hd__nand2_2 _29150_ (.A(_00140_),
    .B(_00313_),
    .Y(_00523_));
 sky130_fd_sc_hd__a211o_2 _29151_ (.A1(_18716_),
    .A2(_00315_),
    .B1(_00314_),
    .C1(_18849_),
    .X(_00524_));
 sky130_fd_sc_hd__and2b_2 _29152_ (.A_N(_00144_),
    .B(_00312_),
    .X(_00525_));
 sky130_fd_sc_hd__and2_2 _29153_ (.A(_00308_),
    .B(_00310_),
    .X(_00527_));
 sky130_fd_sc_hd__nor2_2 _29154_ (.A(_00146_),
    .B(_00311_),
    .Y(_00528_));
 sky130_fd_sc_hd__and2_2 _29155_ (.A(_00149_),
    .B(_00176_),
    .X(_00529_));
 sky130_fd_sc_hd__and2b_2 _29156_ (.A_N(_00147_),
    .B(_00177_),
    .X(_00530_));
 sky130_fd_sc_hd__nor2_2 _29157_ (.A(_00529_),
    .B(_00530_),
    .Y(_00531_));
 sky130_fd_sc_hd__and2b_2 _29158_ (.A_N(_00303_),
    .B(_00305_),
    .X(_00532_));
 sky130_fd_sc_hd__xnor2_2 _29159_ (.A(_00303_),
    .B(_00305_),
    .Y(_00533_));
 sky130_fd_sc_hd__and2_2 _29160_ (.A(_00178_),
    .B(_00533_),
    .X(_00534_));
 sky130_fd_sc_hd__inv_2 _29161_ (.A(_00221_),
    .Y(_00535_));
 sky130_fd_sc_hd__a21o_2 _29162_ (.A1(_00181_),
    .A2(_00535_),
    .B1(_00220_),
    .X(_00536_));
 sky130_fd_sc_hd__nor2_2 _29163_ (.A(_00198_),
    .B(_00199_),
    .Y(_00538_));
 sky130_fd_sc_hd__a21o_2 _29164_ (.A1(_00190_),
    .A2(_00200_),
    .B1(_00538_),
    .X(_00539_));
 sky130_fd_sc_hd__nand2_2 _29165_ (.A(_00152_),
    .B(_00163_),
    .Y(_00540_));
 sky130_fd_sc_hd__o21bai_2 _29166_ (.A1(_00185_),
    .A2(_00187_),
    .B1_N(_00184_),
    .Y(_00541_));
 sky130_fd_sc_hd__or4b_2 _29167_ (.A(_12468_),
    .B(_18120_),
    .C(_18342_),
    .D_N(_18728_),
    .X(_00542_));
 sky130_fd_sc_hd__a22o_2 _29168_ (.A1(_18749_),
    .A2(_18732_),
    .B1(_18728_),
    .B2(_15616_),
    .X(_00543_));
 sky130_fd_sc_hd__a22o_2 _29169_ (.A1(_17392_),
    .A2(_00161_),
    .B1(_00542_),
    .B2(_00543_),
    .X(_00544_));
 sky130_fd_sc_hd__nand4_2 _29170_ (.A(_17392_),
    .B(_00161_),
    .C(_00542_),
    .D(_00543_),
    .Y(_00545_));
 sky130_fd_sc_hd__nand3_2 _29171_ (.A(_00541_),
    .B(_00544_),
    .C(_00545_),
    .Y(_00546_));
 sky130_fd_sc_hd__a21o_2 _29172_ (.A1(_00544_),
    .A2(_00545_),
    .B1(_00541_),
    .X(_00547_));
 sky130_fd_sc_hd__nand3_2 _29173_ (.A(_00540_),
    .B(_00546_),
    .C(_00547_),
    .Y(_00549_));
 sky130_fd_sc_hd__a21o_2 _29174_ (.A1(_00546_),
    .A2(_00547_),
    .B1(_00540_),
    .X(_00550_));
 sky130_fd_sc_hd__nand3_2 _29175_ (.A(_00539_),
    .B(_00549_),
    .C(_00550_),
    .Y(_00551_));
 sky130_fd_sc_hd__a21o_2 _29176_ (.A1(_00549_),
    .A2(_00550_),
    .B1(_00539_),
    .X(_00552_));
 sky130_fd_sc_hd__nand2_2 _29177_ (.A(_00166_),
    .B(_00168_),
    .Y(_00553_));
 sky130_fd_sc_hd__and3_2 _29178_ (.A(_00551_),
    .B(_00552_),
    .C(_00553_),
    .X(_00554_));
 sky130_fd_sc_hd__a21oi_2 _29179_ (.A1(_00551_),
    .A2(_00552_),
    .B1(_00553_),
    .Y(_00555_));
 sky130_fd_sc_hd__o21ba_2 _29180_ (.A1(_18737_),
    .A2(_00171_),
    .B1_N(_00170_),
    .X(_00556_));
 sky130_fd_sc_hd__or3_4 _29181_ (.A(_00554_),
    .B(_00555_),
    .C(_00556_),
    .X(_00557_));
 sky130_fd_sc_hd__o21ai_2 _29182_ (.A1(_00554_),
    .A2(_00555_),
    .B1(_00556_),
    .Y(_00558_));
 sky130_fd_sc_hd__nand2_2 _29183_ (.A(iY[27]),
    .B(iY[59]),
    .Y(_00560_));
 sky130_fd_sc_hd__or2_2 _29184_ (.A(iY[27]),
    .B(iY[59]),
    .X(_00561_));
 sky130_fd_sc_hd__nand2_2 _29185_ (.A(_00560_),
    .B(_00561_),
    .Y(_00562_));
 sky130_fd_sc_hd__o31a_2 _29186_ (.A1(_18724_),
    .A2(_00157_),
    .A3(_00159_),
    .B1(_00155_),
    .X(_00563_));
 sky130_fd_sc_hd__xor2_2 _29187_ (.A(_00562_),
    .B(_00563_),
    .X(_00564_));
 sky130_fd_sc_hd__buf_1 _29188_ (.A(_00564_),
    .X(_00565_));
 sky130_fd_sc_hd__buf_6 _29189_ (.A(_00565_),
    .X(_00566_));
 sky130_fd_sc_hd__buf_6 _29190_ (.A(_00566_),
    .X(_00567_));
 sky130_fd_sc_hd__nand4_2 _29191_ (.A(_14592_),
    .B(_00557_),
    .C(_00558_),
    .D(_00567_),
    .Y(_00568_));
 sky130_fd_sc_hd__a22o_2 _29192_ (.A1(_00557_),
    .A2(_00558_),
    .B1(_00567_),
    .B2(_14592_),
    .X(_00569_));
 sky130_fd_sc_hd__and3_4 _29193_ (.A(_00536_),
    .B(_00568_),
    .C(_00569_),
    .X(_00571_));
 sky130_fd_sc_hd__a21oi_2 _29194_ (.A1(_00568_),
    .A2(_00569_),
    .B1(_00536_),
    .Y(_00572_));
 sky130_fd_sc_hd__and2b_2 _29195_ (.A_N(_00174_),
    .B(_00173_),
    .X(_00573_));
 sky130_fd_sc_hd__nor3b_2 _29196_ (.A(_00571_),
    .B(_00572_),
    .C_N(_00573_),
    .Y(_00574_));
 sky130_fd_sc_hd__o21ba_2 _29197_ (.A1(_00571_),
    .A2(_00572_),
    .B1_N(_00573_),
    .X(_00575_));
 sky130_fd_sc_hd__or2b_2 _29198_ (.A(_00301_),
    .B_N(_00299_),
    .X(_00576_));
 sky130_fd_sc_hd__nand2_2 _29199_ (.A(_00223_),
    .B(_00302_),
    .Y(_00577_));
 sky130_fd_sc_hd__nand2b_2 _29200_ (.A_N(_00225_),
    .B(_00246_),
    .Y(_00578_));
 sky130_fd_sc_hd__and4_2 _29201_ (.A(_15624_),
    .B(_16268_),
    .C(_17629_),
    .D(_18101_),
    .X(_00579_));
 sky130_fd_sc_hd__o22a_2 _29202_ (.A1(_14343_),
    .A2(_17406_),
    .B1(_17627_),
    .B2(_14640_),
    .X(_00580_));
 sky130_fd_sc_hd__or3_4 _29203_ (.A(_14346_),
    .B(_18110_),
    .C(_18112_),
    .X(_00582_));
 sky130_fd_sc_hd__o21a_2 _29204_ (.A1(_00579_),
    .A2(_00580_),
    .B1(_00582_),
    .X(_00583_));
 sky130_fd_sc_hd__or3_4 _29205_ (.A(_00579_),
    .B(_00580_),
    .C(_00582_),
    .X(_00584_));
 sky130_fd_sc_hd__nor2b_2 _29206_ (.A(_00583_),
    .B_N(_00584_),
    .Y(_00585_));
 sky130_fd_sc_hd__or3b_2 _29207_ (.A(_14983_),
    .B(_16616_),
    .C_N(_00192_),
    .X(_00586_));
 sky130_fd_sc_hd__a2bb2o_2 _29208_ (.A1_N(_14983_),
    .A2_N(_16257_),
    .B1(_16613_),
    .B2(_14652_),
    .X(_00587_));
 sky130_fd_sc_hd__nand2_2 _29209_ (.A(_00586_),
    .B(_00587_),
    .Y(_00588_));
 sky130_fd_sc_hd__buf_1 _29210_ (.A(_14357_),
    .X(_00589_));
 sky130_fd_sc_hd__or2_2 _29211_ (.A(_00589_),
    .B(_16922_),
    .X(_00590_));
 sky130_fd_sc_hd__xnor2_2 _29212_ (.A(_00588_),
    .B(_00590_),
    .Y(_00591_));
 sky130_fd_sc_hd__o21a_2 _29213_ (.A1(_00194_),
    .A2(_00196_),
    .B1(_00191_),
    .X(_00593_));
 sky130_fd_sc_hd__xor2_2 _29214_ (.A(_00591_),
    .B(_00593_),
    .X(_00594_));
 sky130_fd_sc_hd__xor2_2 _29215_ (.A(_00585_),
    .B(_00594_),
    .X(_00595_));
 sky130_fd_sc_hd__a2bb2o_2 _29216_ (.A1_N(_00209_),
    .A2_N(_00211_),
    .B1(_18769_),
    .B2(_00207_),
    .X(_00596_));
 sky130_fd_sc_hd__and3_2 _29217_ (.A(_14606_),
    .B(_15679_),
    .C(_18784_),
    .X(_00597_));
 sky130_fd_sc_hd__a21oi_2 _29218_ (.A1(_00231_),
    .A2(_00232_),
    .B1(_00597_),
    .Y(_00598_));
 sky130_fd_sc_hd__nor2_2 _29219_ (.A(_14988_),
    .B(_16237_),
    .Y(_00599_));
 sky130_fd_sc_hd__xnor2_2 _29220_ (.A(_00207_),
    .B(_00599_),
    .Y(_00600_));
 sky130_fd_sc_hd__nor2_2 _29221_ (.A(_15211_),
    .B(_15835_),
    .Y(_00601_));
 sky130_fd_sc_hd__xnor2_2 _29222_ (.A(_00600_),
    .B(_00601_),
    .Y(_00602_));
 sky130_fd_sc_hd__xnor2_2 _29223_ (.A(_00598_),
    .B(_00602_),
    .Y(_00604_));
 sky130_fd_sc_hd__xnor2_2 _29224_ (.A(_00596_),
    .B(_00604_),
    .Y(_00605_));
 sky130_fd_sc_hd__and2_2 _29225_ (.A(_00206_),
    .B(_00212_),
    .X(_00606_));
 sky130_fd_sc_hd__a21oi_2 _29226_ (.A1(_00205_),
    .A2(_00213_),
    .B1(_00606_),
    .Y(_00607_));
 sky130_fd_sc_hd__nor2_2 _29227_ (.A(_00605_),
    .B(_00607_),
    .Y(_00608_));
 sky130_fd_sc_hd__and2_2 _29228_ (.A(_00605_),
    .B(_00607_),
    .X(_00609_));
 sky130_fd_sc_hd__nor2_2 _29229_ (.A(_00608_),
    .B(_00609_),
    .Y(_00610_));
 sky130_fd_sc_hd__and2_2 _29230_ (.A(_00595_),
    .B(_00610_),
    .X(_00611_));
 sky130_fd_sc_hd__nor2_2 _29231_ (.A(_00595_),
    .B(_00610_),
    .Y(_00612_));
 sky130_fd_sc_hd__a211oi_2 _29232_ (.A1(_00244_),
    .A2(_00578_),
    .B1(_00611_),
    .C1(_00612_),
    .Y(_00613_));
 sky130_fd_sc_hd__o211a_2 _29233_ (.A1(_00611_),
    .A2(_00612_),
    .B1(_00244_),
    .C1(_00578_),
    .X(_00615_));
 sky130_fd_sc_hd__a211oi_2 _29234_ (.A1(_00215_),
    .A2(_00217_),
    .B1(_00613_),
    .C1(_00615_),
    .Y(_00616_));
 sky130_fd_sc_hd__o211a_2 _29235_ (.A1(_00613_),
    .A2(_00615_),
    .B1(_00215_),
    .C1(_00217_),
    .X(_00617_));
 sky130_fd_sc_hd__or2_2 _29236_ (.A(_00293_),
    .B(_00297_),
    .X(_00618_));
 sky130_fd_sc_hd__nand2_2 _29237_ (.A(_00247_),
    .B(_00298_),
    .Y(_00619_));
 sky130_fd_sc_hd__or2_2 _29238_ (.A(_00238_),
    .B(_00240_),
    .X(_00620_));
 sky130_fd_sc_hd__o21a_2 _29239_ (.A1(_00233_),
    .A2(_00242_),
    .B1(_00620_),
    .X(_00621_));
 sky130_fd_sc_hd__and2_2 _29240_ (.A(_00249_),
    .B(_00257_),
    .X(_00622_));
 sky130_fd_sc_hd__and3_2 _29241_ (.A(_14608_),
    .B(_17460_),
    .C(_00229_),
    .X(_00623_));
 sky130_fd_sc_hd__and3_2 _29242_ (.A(_14410_),
    .B(_15224_),
    .C(_15226_),
    .X(_00624_));
 sky130_fd_sc_hd__a21oi_2 _29243_ (.A1(_14608_),
    .A2(_15679_),
    .B1(_00624_),
    .Y(_00626_));
 sky130_fd_sc_hd__nor2_2 _29244_ (.A(_00623_),
    .B(_00626_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand2_2 _29245_ (.A(_16292_),
    .B(_15617_),
    .Y(_00628_));
 sky130_fd_sc_hd__xor2_2 _29246_ (.A(_00627_),
    .B(_00628_),
    .X(_00629_));
 sky130_fd_sc_hd__or4_4 _29247_ (.A(_14612_),
    .B(_13893_),
    .C(_17696_),
    .D(_16988_),
    .X(_00630_));
 sky130_fd_sc_hd__a22o_2 _29248_ (.A1(_13888_),
    .A2(_15900_),
    .B1(_17006_),
    .B2(_13543_),
    .X(_00631_));
 sky130_fd_sc_hd__nand2_2 _29249_ (.A(_00630_),
    .B(_00631_),
    .Y(_00632_));
 sky130_fd_sc_hd__buf_1 _29250_ (.A(_15672_),
    .X(_00633_));
 sky130_fd_sc_hd__nand2_2 _29251_ (.A(_14392_),
    .B(_00633_),
    .Y(_00634_));
 sky130_fd_sc_hd__xor2_2 _29252_ (.A(_00632_),
    .B(_00634_),
    .X(_00635_));
 sky130_fd_sc_hd__o21a_2 _29253_ (.A1(_00236_),
    .A2(_00237_),
    .B1(_00234_),
    .X(_00637_));
 sky130_fd_sc_hd__xor2_2 _29254_ (.A(_00635_),
    .B(_00637_),
    .X(_00638_));
 sky130_fd_sc_hd__xor2_2 _29255_ (.A(_00629_),
    .B(_00638_),
    .X(_00639_));
 sky130_fd_sc_hd__o21ai_2 _29256_ (.A1(_00622_),
    .A2(_00259_),
    .B1(_00639_),
    .Y(_00640_));
 sky130_fd_sc_hd__or3_2 _29257_ (.A(_00622_),
    .B(_00259_),
    .C(_00639_),
    .X(_00641_));
 sky130_fd_sc_hd__and2_2 _29258_ (.A(_00640_),
    .B(_00641_),
    .X(_00642_));
 sky130_fd_sc_hd__xnor2_2 _29259_ (.A(_00621_),
    .B(_00642_),
    .Y(_00643_));
 sky130_fd_sc_hd__or2_2 _29260_ (.A(_00289_),
    .B(_00291_),
    .X(_00644_));
 sky130_fd_sc_hd__nand2_2 _29261_ (.A(_00261_),
    .B(_00292_),
    .Y(_00645_));
 sky130_fd_sc_hd__a21bo_2 _29262_ (.A1(_00253_),
    .A2(_00256_),
    .B1_N(_00251_),
    .X(_00646_));
 sky130_fd_sc_hd__a31o_2 _29263_ (.A1(_18192_),
    .A2(_18209_),
    .A3(_00266_),
    .B1(_00264_),
    .X(_00648_));
 sky130_fd_sc_hd__buf_1 _29264_ (.A(_17007_),
    .X(_00649_));
 sky130_fd_sc_hd__nor2_2 _29265_ (.A(_12848_),
    .B(_17482_),
    .Y(_00650_));
 sky130_fd_sc_hd__xnor2_2 _29266_ (.A(_00250_),
    .B(_00650_),
    .Y(_00651_));
 sky130_fd_sc_hd__nor2_2 _29267_ (.A(_00649_),
    .B(_00651_),
    .Y(_00652_));
 sky130_fd_sc_hd__o21a_2 _29268_ (.A1(_14626_),
    .A2(_00649_),
    .B1(_00651_),
    .X(_00653_));
 sky130_fd_sc_hd__a21oi_2 _29269_ (.A1(_17463_),
    .A2(_00652_),
    .B1(_00653_),
    .Y(_00654_));
 sky130_fd_sc_hd__xor2_2 _29270_ (.A(_00648_),
    .B(_00654_),
    .X(_00655_));
 sky130_fd_sc_hd__xor2_2 _29271_ (.A(_00646_),
    .B(_00655_),
    .X(_00656_));
 sky130_fd_sc_hd__nor2_2 _29272_ (.A(_15646_),
    .B(_18443_),
    .Y(_00657_));
 sky130_fd_sc_hd__nor2_2 _29273_ (.A(_15650_),
    .B(_00271_),
    .Y(_00659_));
 sky130_fd_sc_hd__and3_2 _29274_ (.A(_14980_),
    .B(_18203_),
    .C(_00659_),
    .X(_00660_));
 sky130_fd_sc_hd__buf_1 _29275_ (.A(_12243_),
    .X(_00661_));
 sky130_fd_sc_hd__buf_2 _29276_ (.A(_18203_),
    .X(_00662_));
 sky130_fd_sc_hd__a21o_2 _29277_ (.A1(_00661_),
    .A2(_00662_),
    .B1(_00659_),
    .X(_00663_));
 sky130_fd_sc_hd__or2b_2 _29278_ (.A(_00660_),
    .B_N(_00663_),
    .X(_00664_));
 sky130_fd_sc_hd__xnor2_2 _29279_ (.A(_00657_),
    .B(_00664_),
    .Y(_00665_));
 sky130_fd_sc_hd__or2_2 _29280_ (.A(_18822_),
    .B(_18823_),
    .X(_00666_));
 sky130_fd_sc_hd__nor2_2 _29281_ (.A(_11794_),
    .B(_00666_),
    .Y(_00667_));
 sky130_fd_sc_hd__or3_4 _29282_ (.A(_11576_),
    .B(_00278_),
    .C(_00280_),
    .X(_00668_));
 sky130_fd_sc_hd__a311o_2 _29283_ (.A1(_18451_),
    .A2(_18454_),
    .A3(_18819_),
    .B1(_00277_),
    .C1(_18818_),
    .X(_00670_));
 sky130_fd_sc_hd__or2_2 _29284_ (.A(iX[27]),
    .B(iX[59]),
    .X(_00671_));
 sky130_fd_sc_hd__nand2_2 _29285_ (.A(iX[27]),
    .B(iX[59]),
    .Y(_00672_));
 sky130_fd_sc_hd__nand2_2 _29286_ (.A(_00671_),
    .B(_00672_),
    .Y(_00673_));
 sky130_fd_sc_hd__and3_2 _29287_ (.A(_00275_),
    .B(_00670_),
    .C(_00673_),
    .X(_00674_));
 sky130_fd_sc_hd__a21oi_2 _29288_ (.A1(_00275_),
    .A2(_00670_),
    .B1(_00673_),
    .Y(_00675_));
 sky130_fd_sc_hd__or4_4 _29289_ (.A(_11566_),
    .B(_00668_),
    .C(_00674_),
    .D(_00675_),
    .X(_00676_));
 sky130_fd_sc_hd__o31ai_2 _29290_ (.A1(_11567_),
    .A2(_00674_),
    .A3(_00675_),
    .B1(_00668_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand3_2 _29291_ (.A(_00667_),
    .B(_00676_),
    .C(_00677_),
    .Y(_00678_));
 sky130_fd_sc_hd__a21o_2 _29292_ (.A1(_00676_),
    .A2(_00677_),
    .B1(_00667_),
    .X(_00679_));
 sky130_fd_sc_hd__a2bb2o_2 _29293_ (.A1_N(_18824_),
    .A2_N(_00668_),
    .B1(_00282_),
    .B2(_00272_),
    .X(_00681_));
 sky130_fd_sc_hd__nand3_2 _29294_ (.A(_00678_),
    .B(_00679_),
    .C(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__a21o_2 _29295_ (.A1(_00678_),
    .A2(_00679_),
    .B1(_00681_),
    .X(_00683_));
 sky130_fd_sc_hd__nand3_2 _29296_ (.A(_00665_),
    .B(_00682_),
    .C(_00683_),
    .Y(_00684_));
 sky130_fd_sc_hd__a21o_2 _29297_ (.A1(_00682_),
    .A2(_00683_),
    .B1(_00665_),
    .X(_00685_));
 sky130_fd_sc_hd__a21bo_2 _29298_ (.A1(_00267_),
    .A2(_00286_),
    .B1_N(_00284_),
    .X(_00686_));
 sky130_fd_sc_hd__nand3_2 _29299_ (.A(_00684_),
    .B(_00685_),
    .C(_00686_),
    .Y(_00687_));
 sky130_fd_sc_hd__a21o_2 _29300_ (.A1(_00684_),
    .A2(_00685_),
    .B1(_00686_),
    .X(_00688_));
 sky130_fd_sc_hd__and3_2 _29301_ (.A(_00656_),
    .B(_00687_),
    .C(_00688_),
    .X(_00689_));
 sky130_fd_sc_hd__a21oi_2 _29302_ (.A1(_00687_),
    .A2(_00688_),
    .B1(_00656_),
    .Y(_00690_));
 sky130_fd_sc_hd__a211o_2 _29303_ (.A1(_00644_),
    .A2(_00645_),
    .B1(_00689_),
    .C1(_00690_),
    .X(_00692_));
 sky130_fd_sc_hd__o211ai_2 _29304_ (.A1(_00689_),
    .A2(_00690_),
    .B1(_00644_),
    .C1(_00645_),
    .Y(_00693_));
 sky130_fd_sc_hd__and3_2 _29305_ (.A(_00643_),
    .B(_00692_),
    .C(_00693_),
    .X(_00694_));
 sky130_fd_sc_hd__a21oi_2 _29306_ (.A1(_00692_),
    .A2(_00693_),
    .B1(_00643_),
    .Y(_00695_));
 sky130_fd_sc_hd__a211oi_2 _29307_ (.A1(_00618_),
    .A2(_00619_),
    .B1(_00694_),
    .C1(_00695_),
    .Y(_00696_));
 sky130_fd_sc_hd__o211a_2 _29308_ (.A1(_00694_),
    .A2(_00695_),
    .B1(_00618_),
    .C1(_00619_),
    .X(_00697_));
 sky130_fd_sc_hd__nor4_2 _29309_ (.A(_00616_),
    .B(_00617_),
    .C(_00696_),
    .D(_00697_),
    .Y(_00698_));
 sky130_fd_sc_hd__o22a_2 _29310_ (.A1(_00616_),
    .A2(_00617_),
    .B1(_00696_),
    .B2(_00697_),
    .X(_00699_));
 sky130_fd_sc_hd__a211o_2 _29311_ (.A1(_00576_),
    .A2(_00577_),
    .B1(_00698_),
    .C1(_00699_),
    .X(_00700_));
 sky130_fd_sc_hd__o211ai_2 _29312_ (.A1(_00698_),
    .A2(_00699_),
    .B1(_00576_),
    .C1(_00577_),
    .Y(_00701_));
 sky130_fd_sc_hd__nand4bb_2 _29313_ (.A_N(_00574_),
    .B_N(_00575_),
    .C(_00700_),
    .D(_00701_),
    .Y(_00703_));
 sky130_fd_sc_hd__a2bb2o_2 _29314_ (.A1_N(_00574_),
    .A2_N(_00575_),
    .B1(_00700_),
    .B2(_00701_),
    .X(_00704_));
 sky130_fd_sc_hd__o211a_2 _29315_ (.A1(_00532_),
    .A2(_00534_),
    .B1(_00703_),
    .C1(_00704_),
    .X(_00705_));
 sky130_fd_sc_hd__a211oi_2 _29316_ (.A1(_00703_),
    .A2(_00704_),
    .B1(_00532_),
    .C1(_00534_),
    .Y(_00706_));
 sky130_fd_sc_hd__or3_4 _29317_ (.A(_00531_),
    .B(_00705_),
    .C(_00706_),
    .X(_00707_));
 sky130_fd_sc_hd__o21ai_2 _29318_ (.A1(_00705_),
    .A2(_00706_),
    .B1(_00531_),
    .Y(_00708_));
 sky130_fd_sc_hd__o211ai_2 _29319_ (.A1(_00527_),
    .A2(_00528_),
    .B1(_00707_),
    .C1(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__a211o_2 _29320_ (.A1(_00707_),
    .A2(_00708_),
    .B1(_00527_),
    .C1(_00528_),
    .X(_00710_));
 sky130_fd_sc_hd__and3_4 _29321_ (.A(_00525_),
    .B(_00709_),
    .C(_00710_),
    .X(_00711_));
 sky130_fd_sc_hd__a21oi_2 _29322_ (.A1(_00709_),
    .A2(_00710_),
    .B1(_00525_),
    .Y(_00712_));
 sky130_fd_sc_hd__or2_2 _29323_ (.A(_00711_),
    .B(_00712_),
    .X(_00714_));
 sky130_fd_sc_hd__a21o_2 _29324_ (.A1(_00523_),
    .A2(_00524_),
    .B1(_00714_),
    .X(_00715_));
 sky130_fd_sc_hd__nand3_2 _29325_ (.A(_00523_),
    .B(_00524_),
    .C(_00714_),
    .Y(_00716_));
 sky130_fd_sc_hd__inv_2 _29326_ (.A(_00455_),
    .Y(_00717_));
 sky130_fd_sc_hd__nor2_2 _29327_ (.A(_00457_),
    .B(_00458_),
    .Y(_00718_));
 sky130_fd_sc_hd__and3_2 _29328_ (.A(_00430_),
    .B(_00445_),
    .C(_00446_),
    .X(_00719_));
 sky130_fd_sc_hd__inv_2 _29329_ (.A(_00453_),
    .Y(_00720_));
 sky130_fd_sc_hd__or2b_2 _29330_ (.A(_00328_),
    .B_N(_00327_),
    .X(_00721_));
 sky130_fd_sc_hd__and4_2 _29331_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[56]),
    .D(iX[57]),
    .X(_00722_));
 sky130_fd_sc_hd__a22oi_2 _29332_ (.A1(iY[35]),
    .A2(iX[56]),
    .B1(iX[57]),
    .B2(iY[34]),
    .Y(_00723_));
 sky130_fd_sc_hd__nor2_2 _29333_ (.A(_00722_),
    .B(_00723_),
    .Y(_00725_));
 sky130_fd_sc_hd__nand2_2 _29334_ (.A(iY[33]),
    .B(iX[58]),
    .Y(_00726_));
 sky130_fd_sc_hd__xnor2_2 _29335_ (.A(_00725_),
    .B(_00726_),
    .Y(_00727_));
 sky130_fd_sc_hd__o21ba_2 _29336_ (.A1(_00324_),
    .A2(_00326_),
    .B1_N(_00323_),
    .X(_00728_));
 sky130_fd_sc_hd__xnor2_2 _29337_ (.A(_00727_),
    .B(_00728_),
    .Y(_00729_));
 sky130_fd_sc_hd__and2_2 _29338_ (.A(iY[36]),
    .B(iX[59]),
    .X(_00730_));
 sky130_fd_sc_hd__nand3_2 _29339_ (.A(iY[32]),
    .B(iX[55]),
    .C(_00730_),
    .Y(_00731_));
 sky130_fd_sc_hd__a22o_2 _29340_ (.A1(iY[36]),
    .A2(iX[55]),
    .B1(iX[59]),
    .B2(iY[32]),
    .X(_00732_));
 sky130_fd_sc_hd__and2_2 _29341_ (.A(iY[37]),
    .B(iX[54]),
    .X(_00733_));
 sky130_fd_sc_hd__a21oi_2 _29342_ (.A1(_00731_),
    .A2(_00732_),
    .B1(_00733_),
    .Y(_00734_));
 sky130_fd_sc_hd__and3_2 _29343_ (.A(_00731_),
    .B(_00732_),
    .C(_00733_),
    .X(_00736_));
 sky130_fd_sc_hd__nor2_2 _29344_ (.A(_00734_),
    .B(_00736_),
    .Y(_00737_));
 sky130_fd_sc_hd__xnor2_2 _29345_ (.A(_00729_),
    .B(_00737_),
    .Y(_00738_));
 sky130_fd_sc_hd__a21o_2 _29346_ (.A1(_00721_),
    .A2(_00336_),
    .B1(_00738_),
    .X(_00739_));
 sky130_fd_sc_hd__nand3_2 _29347_ (.A(_00721_),
    .B(_00336_),
    .C(_00738_),
    .Y(_00740_));
 sky130_fd_sc_hd__o21ba_2 _29348_ (.A1(_00345_),
    .A2(_00347_),
    .B1_N(_00344_),
    .X(_00741_));
 sky130_fd_sc_hd__o21ba_2 _29349_ (.A1(_00332_),
    .A2(_00334_),
    .B1_N(_00331_),
    .X(_00742_));
 sky130_fd_sc_hd__and4_2 _29350_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[52]),
    .D(iX[53]),
    .X(_00743_));
 sky130_fd_sc_hd__a22oi_2 _29351_ (.A1(iY[39]),
    .A2(iX[52]),
    .B1(iX[53]),
    .B2(iY[38]),
    .Y(_00744_));
 sky130_fd_sc_hd__nor2_2 _29352_ (.A(_00743_),
    .B(_00744_),
    .Y(_00745_));
 sky130_fd_sc_hd__nand2_2 _29353_ (.A(iY[40]),
    .B(iX[51]),
    .Y(_00747_));
 sky130_fd_sc_hd__xnor2_2 _29354_ (.A(_00745_),
    .B(_00747_),
    .Y(_00748_));
 sky130_fd_sc_hd__xnor2_2 _29355_ (.A(_00742_),
    .B(_00748_),
    .Y(_00749_));
 sky130_fd_sc_hd__xnor2_2 _29356_ (.A(_00741_),
    .B(_00749_),
    .Y(_00750_));
 sky130_fd_sc_hd__nand3_2 _29357_ (.A(_00739_),
    .B(_00740_),
    .C(_00750_),
    .Y(_00751_));
 sky130_fd_sc_hd__a21o_2 _29358_ (.A1(_00739_),
    .A2(_00740_),
    .B1(_00750_),
    .X(_00752_));
 sky130_fd_sc_hd__nand2_2 _29359_ (.A(_00751_),
    .B(_00752_),
    .Y(_00753_));
 sky130_fd_sc_hd__a21bo_2 _29360_ (.A1(_00341_),
    .A2(_00350_),
    .B1_N(_00339_),
    .X(_00754_));
 sky130_fd_sc_hd__xor2_2 _29361_ (.A(_00753_),
    .B(_00754_),
    .X(_00755_));
 sky130_fd_sc_hd__a21bo_2 _29362_ (.A1(_00365_),
    .A2(_00374_),
    .B1_N(_00371_),
    .X(_00756_));
 sky130_fd_sc_hd__or2b_2 _29363_ (.A(_00343_),
    .B_N(_00348_),
    .X(_00758_));
 sky130_fd_sc_hd__or2b_2 _29364_ (.A(_00342_),
    .B_N(_00349_),
    .X(_00759_));
 sky130_fd_sc_hd__and4_2 _29365_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[46]),
    .D(iX[47]),
    .X(_00760_));
 sky130_fd_sc_hd__a22oi_2 _29366_ (.A1(iY[45]),
    .A2(iX[46]),
    .B1(iX[47]),
    .B2(iY[44]),
    .Y(_00761_));
 sky130_fd_sc_hd__nor2_2 _29367_ (.A(_00760_),
    .B(_00761_),
    .Y(_00762_));
 sky130_fd_sc_hd__nand2_2 _29368_ (.A(iX[45]),
    .B(iY[46]),
    .Y(_00763_));
 sky130_fd_sc_hd__xnor2_2 _29369_ (.A(_00762_),
    .B(_00763_),
    .Y(_00764_));
 sky130_fd_sc_hd__and4_2 _29370_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[49]),
    .D(iX[50]),
    .X(_00765_));
 sky130_fd_sc_hd__a22oi_2 _29371_ (.A1(iY[42]),
    .A2(iX[49]),
    .B1(iX[50]),
    .B2(iY[41]),
    .Y(_00766_));
 sky130_fd_sc_hd__nor2_2 _29372_ (.A(_00765_),
    .B(_00766_),
    .Y(_00767_));
 sky130_fd_sc_hd__nand2_2 _29373_ (.A(iY[43]),
    .B(iX[48]),
    .Y(_00769_));
 sky130_fd_sc_hd__xnor2_2 _29374_ (.A(_00767_),
    .B(_00769_),
    .Y(_00770_));
 sky130_fd_sc_hd__o21ba_2 _29375_ (.A1(_00367_),
    .A2(_00369_),
    .B1_N(_00366_),
    .X(_00771_));
 sky130_fd_sc_hd__xnor2_2 _29376_ (.A(_00770_),
    .B(_00771_),
    .Y(_00772_));
 sky130_fd_sc_hd__and2_2 _29377_ (.A(_00764_),
    .B(_00772_),
    .X(_00773_));
 sky130_fd_sc_hd__nor2_2 _29378_ (.A(_00764_),
    .B(_00772_),
    .Y(_00774_));
 sky130_fd_sc_hd__or2_2 _29379_ (.A(_00773_),
    .B(_00774_),
    .X(_00775_));
 sky130_fd_sc_hd__a21o_2 _29380_ (.A1(_00758_),
    .A2(_00759_),
    .B1(_00775_),
    .X(_00776_));
 sky130_fd_sc_hd__and3_2 _29381_ (.A(_00758_),
    .B(_00759_),
    .C(_00775_),
    .X(_00777_));
 sky130_fd_sc_hd__inv_2 _29382_ (.A(_00777_),
    .Y(_00778_));
 sky130_fd_sc_hd__nand3_2 _29383_ (.A(_00756_),
    .B(_00776_),
    .C(_00778_),
    .Y(_00780_));
 sky130_fd_sc_hd__a21o_2 _29384_ (.A1(_00776_),
    .A2(_00778_),
    .B1(_00756_),
    .X(_00781_));
 sky130_fd_sc_hd__nand2_2 _29385_ (.A(_00780_),
    .B(_00781_),
    .Y(_00782_));
 sky130_fd_sc_hd__nor2_2 _29386_ (.A(_00755_),
    .B(_00782_),
    .Y(_00783_));
 sky130_fd_sc_hd__and2_2 _29387_ (.A(_00755_),
    .B(_00782_),
    .X(_00784_));
 sky130_fd_sc_hd__nor2_2 _29388_ (.A(_00783_),
    .B(_00784_),
    .Y(_00785_));
 sky130_fd_sc_hd__a21bo_2 _29389_ (.A1(_00354_),
    .A2(_00355_),
    .B1_N(_00381_),
    .X(_00786_));
 sky130_fd_sc_hd__xnor2_2 _29390_ (.A(_00785_),
    .B(_00786_),
    .Y(_00787_));
 sky130_fd_sc_hd__and4_2 _29391_ (.A(iX[37]),
    .B(iX[38]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_00788_));
 sky130_fd_sc_hd__a22oi_2 _29392_ (.A1(iX[38]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[37]),
    .Y(_00789_));
 sky130_fd_sc_hd__nor2_2 _29393_ (.A(_00788_),
    .B(_00789_),
    .Y(_00791_));
 sky130_fd_sc_hd__nand2_2 _29394_ (.A(iX[36]),
    .B(iY[55]),
    .Y(_00792_));
 sky130_fd_sc_hd__xnor2_2 _29395_ (.A(_00791_),
    .B(_00792_),
    .Y(_00793_));
 sky130_fd_sc_hd__and4_2 _29396_ (.A(iX[40]),
    .B(iX[41]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_00794_));
 sky130_fd_sc_hd__a22oi_2 _29397_ (.A1(iX[41]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[40]),
    .Y(_00795_));
 sky130_fd_sc_hd__nor2_2 _29398_ (.A(_00794_),
    .B(_00795_),
    .Y(_00796_));
 sky130_fd_sc_hd__nand2_2 _29399_ (.A(iX[39]),
    .B(iY[52]),
    .Y(_00797_));
 sky130_fd_sc_hd__xnor2_2 _29400_ (.A(_00796_),
    .B(_00797_),
    .Y(_00798_));
 sky130_fd_sc_hd__o21ba_2 _29401_ (.A1(_00394_),
    .A2(_00397_),
    .B1_N(_00393_),
    .X(_00799_));
 sky130_fd_sc_hd__xnor2_2 _29402_ (.A(_00798_),
    .B(_00799_),
    .Y(_00800_));
 sky130_fd_sc_hd__and2_2 _29403_ (.A(_00793_),
    .B(_00800_),
    .X(_00802_));
 sky130_fd_sc_hd__nor2_2 _29404_ (.A(_00793_),
    .B(_00800_),
    .Y(_00803_));
 sky130_fd_sc_hd__or2_2 _29405_ (.A(_00802_),
    .B(_00803_),
    .X(_00804_));
 sky130_fd_sc_hd__or3_2 _29406_ (.A(_00405_),
    .B(_00409_),
    .C(_00410_),
    .X(_00805_));
 sky130_fd_sc_hd__o21ba_2 _29407_ (.A1(_00361_),
    .A2(_00364_),
    .B1_N(_00360_),
    .X(_00806_));
 sky130_fd_sc_hd__and4_2 _29408_ (.A(iX[43]),
    .B(iX[44]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_00807_));
 sky130_fd_sc_hd__a22oi_2 _29409_ (.A1(iX[44]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[43]),
    .Y(_00808_));
 sky130_fd_sc_hd__and4bb_2 _29410_ (.A_N(_00807_),
    .B_N(_00808_),
    .C(iX[42]),
    .D(iY[49]),
    .X(_00809_));
 sky130_fd_sc_hd__o2bb2a_2 _29411_ (.A1_N(iX[42]),
    .A2_N(iY[49]),
    .B1(_00807_),
    .B2(_00808_),
    .X(_00810_));
 sky130_fd_sc_hd__nor2_2 _29412_ (.A(_00809_),
    .B(_00810_),
    .Y(_00811_));
 sky130_fd_sc_hd__xnor2_2 _29413_ (.A(_00806_),
    .B(_00811_),
    .Y(_00813_));
 sky130_fd_sc_hd__o21ai_2 _29414_ (.A1(_00407_),
    .A2(_00409_),
    .B1(_00813_),
    .Y(_00814_));
 sky130_fd_sc_hd__or3_2 _29415_ (.A(_00407_),
    .B(_00409_),
    .C(_00813_),
    .X(_00815_));
 sky130_fd_sc_hd__nand2_2 _29416_ (.A(_00814_),
    .B(_00815_),
    .Y(_00816_));
 sky130_fd_sc_hd__a21oi_2 _29417_ (.A1(_00805_),
    .A2(_00413_),
    .B1(_00816_),
    .Y(_00817_));
 sky130_fd_sc_hd__and3_2 _29418_ (.A(_00805_),
    .B(_00413_),
    .C(_00816_),
    .X(_00818_));
 sky130_fd_sc_hd__or3_2 _29419_ (.A(_00804_),
    .B(_00817_),
    .C(_00818_),
    .X(_00819_));
 sky130_fd_sc_hd__o21ai_2 _29420_ (.A1(_00817_),
    .A2(_00818_),
    .B1(_00804_),
    .Y(_00820_));
 sky130_fd_sc_hd__o211a_2 _29421_ (.A1(_00376_),
    .A2(_00379_),
    .B1(_00819_),
    .C1(_00820_),
    .X(_00821_));
 sky130_fd_sc_hd__inv_2 _29422_ (.A(_00821_),
    .Y(_00822_));
 sky130_fd_sc_hd__a211o_2 _29423_ (.A1(_00819_),
    .A2(_00820_),
    .B1(_00376_),
    .C1(_00379_),
    .X(_00824_));
 sky130_fd_sc_hd__o211a_2 _29424_ (.A1(_00416_),
    .A2(_00419_),
    .B1(_00822_),
    .C1(_00824_),
    .X(_00825_));
 sky130_fd_sc_hd__a211oi_2 _29425_ (.A1(_00822_),
    .A2(_00824_),
    .B1(_00416_),
    .C1(_00419_),
    .Y(_00826_));
 sky130_fd_sc_hd__or3_2 _29426_ (.A(_00787_),
    .B(_00825_),
    .C(_00826_),
    .X(_00827_));
 sky130_fd_sc_hd__o21ai_2 _29427_ (.A1(_00825_),
    .A2(_00826_),
    .B1(_00787_),
    .Y(_00828_));
 sky130_fd_sc_hd__and2_2 _29428_ (.A(_00827_),
    .B(_00828_),
    .X(_00829_));
 sky130_fd_sc_hd__o21ai_2 _29429_ (.A1(_00385_),
    .A2(_00425_),
    .B1(_00829_),
    .Y(_00830_));
 sky130_fd_sc_hd__or3_2 _29430_ (.A(_00385_),
    .B(_00425_),
    .C(_00829_),
    .X(_00831_));
 sky130_fd_sc_hd__and2b_2 _29431_ (.A_N(_00399_),
    .B(_00398_),
    .X(_00832_));
 sky130_fd_sc_hd__o21ba_2 _29432_ (.A1(_00434_),
    .A2(_00436_),
    .B1_N(_00433_),
    .X(_00833_));
 sky130_fd_sc_hd__o21ba_2 _29433_ (.A1(_00389_),
    .A2(_00391_),
    .B1_N(_00388_),
    .X(_00835_));
 sky130_fd_sc_hd__and4_2 _29434_ (.A(iX[34]),
    .B(iX[35]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_00836_));
 sky130_fd_sc_hd__a22oi_2 _29435_ (.A1(iX[35]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[34]),
    .Y(_00837_));
 sky130_fd_sc_hd__nor2_2 _29436_ (.A(_00836_),
    .B(_00837_),
    .Y(_00838_));
 sky130_fd_sc_hd__nand2_2 _29437_ (.A(iX[33]),
    .B(iY[58]),
    .Y(_00839_));
 sky130_fd_sc_hd__xnor2_2 _29438_ (.A(_00838_),
    .B(_00839_),
    .Y(_00840_));
 sky130_fd_sc_hd__xnor2_2 _29439_ (.A(_00835_),
    .B(_00840_),
    .Y(_00841_));
 sky130_fd_sc_hd__xnor2_2 _29440_ (.A(_00833_),
    .B(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__o21a_2 _29441_ (.A1(_00832_),
    .A2(_00401_),
    .B1(_00842_),
    .X(_00843_));
 sky130_fd_sc_hd__nor3_2 _29442_ (.A(_00832_),
    .B(_00401_),
    .C(_00842_),
    .Y(_00844_));
 sky130_fd_sc_hd__and2b_2 _29443_ (.A_N(_00432_),
    .B(_00437_),
    .X(_00846_));
 sky130_fd_sc_hd__a21oi_2 _29444_ (.A1(_00042_),
    .A2(_00438_),
    .B1(_00846_),
    .Y(_00847_));
 sky130_fd_sc_hd__nor3_2 _29445_ (.A(_00843_),
    .B(_00844_),
    .C(_00847_),
    .Y(_00848_));
 sky130_fd_sc_hd__o21a_2 _29446_ (.A1(_00843_),
    .A2(_00844_),
    .B1(_00847_),
    .X(_00849_));
 sky130_fd_sc_hd__or2_2 _29447_ (.A(_00848_),
    .B(_00849_),
    .X(_00850_));
 sky130_fd_sc_hd__a21oi_2 _29448_ (.A1(_00045_),
    .A2(_00443_),
    .B1(_00441_),
    .Y(_00851_));
 sky130_fd_sc_hd__or2_2 _29449_ (.A(_00850_),
    .B(_00851_),
    .X(_00852_));
 sky130_fd_sc_hd__nand2_2 _29450_ (.A(_00850_),
    .B(_00851_),
    .Y(_00853_));
 sky130_fd_sc_hd__nand2_2 _29451_ (.A(_00852_),
    .B(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hd__nand2_2 _29452_ (.A(iX[32]),
    .B(iY[59]),
    .Y(_00855_));
 sky130_fd_sc_hd__or2_2 _29453_ (.A(_00854_),
    .B(_00855_),
    .X(_00857_));
 sky130_fd_sc_hd__nand2_2 _29454_ (.A(_00854_),
    .B(_00855_),
    .Y(_00858_));
 sky130_fd_sc_hd__and2_2 _29455_ (.A(_00857_),
    .B(_00858_),
    .X(_00859_));
 sky130_fd_sc_hd__o21a_2 _29456_ (.A1(_00421_),
    .A2(_00423_),
    .B1(_00859_),
    .X(_00860_));
 sky130_fd_sc_hd__nor3_2 _29457_ (.A(_00421_),
    .B(_00423_),
    .C(_00859_),
    .Y(_00861_));
 sky130_fd_sc_hd__o21ai_2 _29458_ (.A1(_00860_),
    .A2(_00861_),
    .B1(_00445_),
    .Y(_00862_));
 sky130_fd_sc_hd__or3_2 _29459_ (.A(_00445_),
    .B(_00860_),
    .C(_00861_),
    .X(_00863_));
 sky130_fd_sc_hd__nand4_2 _29460_ (.A(_00830_),
    .B(_00831_),
    .C(_00862_),
    .D(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__a22o_2 _29461_ (.A1(_00830_),
    .A2(_00831_),
    .B1(_00862_),
    .B2(_00863_),
    .X(_00865_));
 sky130_fd_sc_hd__o211ai_2 _29462_ (.A1(_00427_),
    .A2(_00720_),
    .B1(_00864_),
    .C1(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__a211o_2 _29463_ (.A1(_00864_),
    .A2(_00865_),
    .B1(_00427_),
    .C1(_00720_),
    .X(_00868_));
 sky130_fd_sc_hd__o211ai_2 _29464_ (.A1(_00719_),
    .A2(_00451_),
    .B1(_00866_),
    .C1(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__a211o_2 _29465_ (.A1(_00866_),
    .A2(_00868_),
    .B1(_00719_),
    .C1(_00451_),
    .X(_00870_));
 sky130_fd_sc_hd__o211ai_2 _29466_ (.A1(_00717_),
    .A2(_00718_),
    .B1(_00869_),
    .C1(_00870_),
    .Y(_00871_));
 sky130_fd_sc_hd__a211o_2 _29467_ (.A1(_00869_),
    .A2(_00870_),
    .B1(_00717_),
    .C1(_00718_),
    .X(_00872_));
 sky130_fd_sc_hd__a21oi_2 _29468_ (.A1(_00871_),
    .A2(_00872_),
    .B1(_00460_),
    .Y(_00873_));
 sky130_fd_sc_hd__inv_2 _29469_ (.A(_00464_),
    .Y(_00874_));
 sky130_fd_sc_hd__or3_2 _29470_ (.A(_00070_),
    .B(_00460_),
    .C(_00462_),
    .X(_00875_));
 sky130_fd_sc_hd__o21a_2 _29471_ (.A1(_00874_),
    .A2(_00468_),
    .B1(_00875_),
    .X(_00876_));
 sky130_fd_sc_hd__and3_2 _29472_ (.A(_00460_),
    .B(_00871_),
    .C(_00872_),
    .X(_00877_));
 sky130_fd_sc_hd__nor2_2 _29473_ (.A(_00877_),
    .B(_00873_),
    .Y(_00879_));
 sky130_fd_sc_hd__inv_2 _29474_ (.A(_00879_),
    .Y(_00880_));
 sky130_fd_sc_hd__nand2_2 _29475_ (.A(_00880_),
    .B(_00876_),
    .Y(_00881_));
 sky130_fd_sc_hd__o21ai_2 _29476_ (.A1(_00873_),
    .A2(_00876_),
    .B1(_00881_),
    .Y(_00882_));
 sky130_fd_sc_hd__a21oi_2 _29477_ (.A1(_00715_),
    .A2(_00716_),
    .B1(_00882_),
    .Y(_00883_));
 sky130_fd_sc_hd__and3_2 _29478_ (.A(_00715_),
    .B(_00716_),
    .C(_00882_),
    .X(_00884_));
 sky130_fd_sc_hd__or3_2 _29479_ (.A(oO[27]),
    .B(_00883_),
    .C(_00884_),
    .X(_00885_));
 sky130_fd_sc_hd__o21ai_2 _29480_ (.A1(_00883_),
    .A2(_00884_),
    .B1(oO[27]),
    .Y(_00886_));
 sky130_fd_sc_hd__nor2_2 _29481_ (.A(_00317_),
    .B(_00469_),
    .Y(_00887_));
 sky130_fd_sc_hd__a21o_2 _29482_ (.A1(_10382_),
    .A2(_00470_),
    .B1(_00887_),
    .X(_00888_));
 sky130_fd_sc_hd__a21o_2 _29483_ (.A1(_00885_),
    .A2(_00886_),
    .B1(_00888_),
    .X(_00890_));
 sky130_fd_sc_hd__and3_2 _29484_ (.A(_00885_),
    .B(_00886_),
    .C(_00888_),
    .X(_00891_));
 sky130_fd_sc_hd__inv_2 _29485_ (.A(_00891_),
    .Y(_00892_));
 sky130_fd_sc_hd__nand2_2 _29486_ (.A(_00890_),
    .B(_00892_),
    .Y(_00893_));
 sky130_fd_sc_hd__a21oi_2 _29487_ (.A1(_00474_),
    .A2(_00480_),
    .B1(_00473_),
    .Y(_00894_));
 sky130_fd_sc_hd__xnor2_2 _29488_ (.A(_00893_),
    .B(_00894_),
    .Y(_00895_));
 sky130_fd_sc_hd__xor2_2 _29489_ (.A(_00522_),
    .B(_00895_),
    .X(_00896_));
 sky130_fd_sc_hd__nor2_2 _29490_ (.A(_00482_),
    .B(_00486_),
    .Y(_00897_));
 sky130_fd_sc_hd__xnor2_2 _29491_ (.A(_00896_),
    .B(_00897_),
    .Y(oO[59]));
 sky130_fd_sc_hd__or2b_2 _29492_ (.A(_00514_),
    .B_N(_00516_),
    .X(_00898_));
 sky130_fd_sc_hd__inv_2 _29493_ (.A(_00509_),
    .Y(_00900_));
 sky130_fd_sc_hd__and3_2 _29494_ (.A(iY[29]),
    .B(iX[31]),
    .C(_00103_),
    .X(_00901_));
 sky130_fd_sc_hd__nand2_2 _29495_ (.A(iX[30]),
    .B(iY[30]),
    .Y(_00902_));
 sky130_fd_sc_hd__xor2_2 _29496_ (.A(_00901_),
    .B(_00902_),
    .X(_00903_));
 sky130_fd_sc_hd__o21ba_2 _29497_ (.A1(_00496_),
    .A2(_00498_),
    .B1_N(_00495_),
    .X(_00904_));
 sky130_fd_sc_hd__xnor2_2 _29498_ (.A(_00903_),
    .B(_00904_),
    .Y(_00905_));
 sky130_fd_sc_hd__nand2_2 _29499_ (.A(iX[29]),
    .B(iY[31]),
    .Y(_00906_));
 sky130_fd_sc_hd__and2_2 _29500_ (.A(_00905_),
    .B(_00906_),
    .X(_00907_));
 sky130_fd_sc_hd__nor2_2 _29501_ (.A(_00905_),
    .B(_00906_),
    .Y(_00908_));
 sky130_fd_sc_hd__nor2_2 _29502_ (.A(_00907_),
    .B(_00908_),
    .Y(_00909_));
 sky130_fd_sc_hd__nand2_2 _29503_ (.A(_00510_),
    .B(_00909_),
    .Y(_00911_));
 sky130_fd_sc_hd__or2_2 _29504_ (.A(_00510_),
    .B(_00909_),
    .X(_00912_));
 sky130_fd_sc_hd__nand2_2 _29505_ (.A(_00911_),
    .B(_00912_),
    .Y(_00913_));
 sky130_fd_sc_hd__nor2_2 _29506_ (.A(_00900_),
    .B(_00913_),
    .Y(_00914_));
 sky130_fd_sc_hd__and2_2 _29507_ (.A(_00900_),
    .B(_00913_),
    .X(_00915_));
 sky130_fd_sc_hd__nor2_2 _29508_ (.A(_00914_),
    .B(_00915_),
    .Y(_00916_));
 sky130_fd_sc_hd__o21ba_2 _29509_ (.A1(_00499_),
    .A2(_00501_),
    .B1_N(_00506_),
    .X(_00917_));
 sky130_fd_sc_hd__xor2_2 _29510_ (.A(_00916_),
    .B(_00917_),
    .X(_00918_));
 sky130_fd_sc_hd__a21oi_2 _29511_ (.A1(_00512_),
    .A2(_00898_),
    .B1(_00918_),
    .Y(_00919_));
 sky130_fd_sc_hd__and3_2 _29512_ (.A(_00512_),
    .B(_00898_),
    .C(_00918_),
    .X(_00920_));
 sky130_fd_sc_hd__or2_2 _29513_ (.A(_00919_),
    .B(_00920_),
    .X(_00921_));
 sky130_fd_sc_hd__inv_2 _29514_ (.A(_00519_),
    .Y(_00922_));
 sky130_fd_sc_hd__o31a_2 _29515_ (.A1(_00133_),
    .A2(_00136_),
    .A3(_00518_),
    .B1(_00922_),
    .X(_00923_));
 sky130_fd_sc_hd__xnor2_2 _29516_ (.A(_00921_),
    .B(_00923_),
    .Y(_00924_));
 sky130_fd_sc_hd__nor2_2 _29517_ (.A(_00473_),
    .B(_00891_),
    .Y(_00925_));
 sky130_fd_sc_hd__a21oi_2 _29518_ (.A1(_00474_),
    .A2(_00890_),
    .B1(_00891_),
    .Y(_00926_));
 sky130_fd_sc_hd__a31oi_2 _29519_ (.A1(_00477_),
    .A2(_00479_),
    .A3(_00925_),
    .B1(_00926_),
    .Y(_00927_));
 sky130_fd_sc_hd__nor3_2 _29520_ (.A(_00531_),
    .B(_00705_),
    .C(_00706_),
    .Y(_00928_));
 sky130_fd_sc_hd__nor2_2 _29521_ (.A(iY[27]),
    .B(iY[59]),
    .Y(_00929_));
 sky130_fd_sc_hd__or2_2 _29522_ (.A(_00157_),
    .B(_00562_),
    .X(_00930_));
 sky130_fd_sc_hd__or3_2 _29523_ (.A(_18724_),
    .B(_00158_),
    .C(_00930_),
    .X(_00932_));
 sky130_fd_sc_hd__o211a_2 _29524_ (.A1(_00155_),
    .A2(_00929_),
    .B1(_00932_),
    .C1(_00560_),
    .X(_00933_));
 sky130_fd_sc_hd__a2111o_2 _29525_ (.A1(_16912_),
    .A2(_16916_),
    .B1(_16920_),
    .C1(_17403_),
    .D1(_18334_),
    .X(_00934_));
 sky130_fd_sc_hd__or3_2 _29526_ (.A(_18333_),
    .B(_18726_),
    .C(_00930_),
    .X(_00935_));
 sky130_fd_sc_hd__a21o_2 _29527_ (.A1(_18336_),
    .A2(_00934_),
    .B1(_00935_),
    .X(_00936_));
 sky130_fd_sc_hd__and2_2 _29528_ (.A(iY[28]),
    .B(iY[60]),
    .X(_00937_));
 sky130_fd_sc_hd__nor2_2 _29529_ (.A(iY[28]),
    .B(iY[60]),
    .Y(_00938_));
 sky130_fd_sc_hd__or2_2 _29530_ (.A(_00937_),
    .B(_00938_),
    .X(_00939_));
 sky130_fd_sc_hd__a21oi_2 _29531_ (.A1(_00933_),
    .A2(_00936_),
    .B1(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__and3_2 _29532_ (.A(_00939_),
    .B(_00933_),
    .C(_00936_),
    .X(_00941_));
 sky130_fd_sc_hd__or2_4 _29533_ (.A(_00940_),
    .B(_00941_),
    .X(_00943_));
 sky130_fd_sc_hd__buf_1 _29534_ (.A(_00943_),
    .X(_00944_));
 sky130_fd_sc_hd__nand2_2 _29535_ (.A(_17392_),
    .B(_00566_),
    .Y(_00945_));
 sky130_fd_sc_hd__o21ai_2 _29536_ (.A1(_11579_),
    .A2(_00944_),
    .B1(_00945_),
    .Y(_00946_));
 sky130_fd_sc_hd__or3_2 _29537_ (.A(_11579_),
    .B(_00945_),
    .C(_00943_),
    .X(_00947_));
 sky130_fd_sc_hd__nand2_2 _29538_ (.A(_00946_),
    .B(_00947_),
    .Y(_00948_));
 sky130_fd_sc_hd__nand3_2 _29539_ (.A(_00551_),
    .B(_00552_),
    .C(_00553_),
    .Y(_00949_));
 sky130_fd_sc_hd__nand2_2 _29540_ (.A(_00546_),
    .B(_00549_),
    .Y(_00950_));
 sky130_fd_sc_hd__nor2_2 _29541_ (.A(_00591_),
    .B(_00593_),
    .Y(_00951_));
 sky130_fd_sc_hd__a21o_2 _29542_ (.A1(_00585_),
    .A2(_00594_),
    .B1(_00951_),
    .X(_00952_));
 sky130_fd_sc_hd__nand2_2 _29543_ (.A(_00542_),
    .B(_00545_),
    .Y(_00954_));
 sky130_fd_sc_hd__o21bai_2 _29544_ (.A1(_00580_),
    .A2(_00582_),
    .B1_N(_00579_),
    .Y(_00955_));
 sky130_fd_sc_hd__or4b_2 _29545_ (.A(_15167_),
    .B(_14346_),
    .C(_18342_),
    .D_N(_18728_),
    .X(_00956_));
 sky130_fd_sc_hd__a22o_2 _29546_ (.A1(_14628_),
    .A2(_18732_),
    .B1(_18728_),
    .B2(_18749_),
    .X(_00957_));
 sky130_fd_sc_hd__a22o_2 _29547_ (.A1(_15616_),
    .A2(_00161_),
    .B1(_00956_),
    .B2(_00957_),
    .X(_00958_));
 sky130_fd_sc_hd__nand4_2 _29548_ (.A(_15616_),
    .B(_00161_),
    .C(_00956_),
    .D(_00957_),
    .Y(_00959_));
 sky130_fd_sc_hd__nand3_2 _29549_ (.A(_00955_),
    .B(_00958_),
    .C(_00959_),
    .Y(_00960_));
 sky130_fd_sc_hd__a21o_2 _29550_ (.A1(_00958_),
    .A2(_00959_),
    .B1(_00955_),
    .X(_00961_));
 sky130_fd_sc_hd__nand3_2 _29551_ (.A(_00954_),
    .B(_00960_),
    .C(_00961_),
    .Y(_00962_));
 sky130_fd_sc_hd__a21o_2 _29552_ (.A1(_00960_),
    .A2(_00961_),
    .B1(_00954_),
    .X(_00963_));
 sky130_fd_sc_hd__nand3_2 _29553_ (.A(_00952_),
    .B(_00962_),
    .C(_00963_),
    .Y(_00965_));
 sky130_fd_sc_hd__a21o_2 _29554_ (.A1(_00962_),
    .A2(_00963_),
    .B1(_00952_),
    .X(_00966_));
 sky130_fd_sc_hd__and3_2 _29555_ (.A(_00950_),
    .B(_00965_),
    .C(_00966_),
    .X(_00967_));
 sky130_fd_sc_hd__a21oi_2 _29556_ (.A1(_00965_),
    .A2(_00966_),
    .B1(_00950_),
    .Y(_00968_));
 sky130_fd_sc_hd__a211oi_2 _29557_ (.A1(_00551_),
    .A2(_00949_),
    .B1(_00967_),
    .C1(_00968_),
    .Y(_00969_));
 sky130_fd_sc_hd__o211a_2 _29558_ (.A1(_00967_),
    .A2(_00968_),
    .B1(_00551_),
    .C1(_00949_),
    .X(_00970_));
 sky130_fd_sc_hd__or3_4 _29559_ (.A(_00948_),
    .B(_00969_),
    .C(_00970_),
    .X(_00971_));
 sky130_fd_sc_hd__o21ai_2 _29560_ (.A1(_00969_),
    .A2(_00970_),
    .B1(_00948_),
    .Y(_00972_));
 sky130_fd_sc_hd__o211a_2 _29561_ (.A1(_00613_),
    .A2(_00616_),
    .B1(_00971_),
    .C1(_00972_),
    .X(_00973_));
 sky130_fd_sc_hd__a211oi_2 _29562_ (.A1(_00971_),
    .A2(_00972_),
    .B1(_00613_),
    .C1(_00616_),
    .Y(_00974_));
 sky130_fd_sc_hd__a211o_2 _29563_ (.A1(_00557_),
    .A2(_00568_),
    .B1(_00973_),
    .C1(_00974_),
    .X(_00976_));
 sky130_fd_sc_hd__o211ai_2 _29564_ (.A1(_00973_),
    .A2(_00974_),
    .B1(_00557_),
    .C1(_00568_),
    .Y(_00977_));
 sky130_fd_sc_hd__or2b_2 _29565_ (.A(_00621_),
    .B_N(_00642_),
    .X(_00978_));
 sky130_fd_sc_hd__and4_2 _29566_ (.A(_16268_),
    .B(_16277_),
    .C(_17630_),
    .D(_18101_),
    .X(_00979_));
 sky130_fd_sc_hd__o22a_2 _29567_ (.A1(_00589_),
    .A2(_17408_),
    .B1(_17627_),
    .B2(_00195_),
    .X(_00980_));
 sky130_fd_sc_hd__or3_4 _29568_ (.A(_14640_),
    .B(_18110_),
    .C(_18112_),
    .X(_00981_));
 sky130_fd_sc_hd__o21a_2 _29569_ (.A1(_00979_),
    .A2(_00980_),
    .B1(_00981_),
    .X(_00982_));
 sky130_fd_sc_hd__or3_4 _29570_ (.A(_00979_),
    .B(_00980_),
    .C(_00981_),
    .X(_00983_));
 sky130_fd_sc_hd__nor2b_2 _29571_ (.A(_00982_),
    .B_N(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hd__nor2_2 _29572_ (.A(_15211_),
    .B(_16255_),
    .Y(_00985_));
 sky130_fd_sc_hd__or3b_2 _29573_ (.A(_14983_),
    .B(_16617_),
    .C_N(_00985_),
    .X(_00987_));
 sky130_fd_sc_hd__a21o_2 _29574_ (.A1(_14648_),
    .A2(_16613_),
    .B1(_00985_),
    .X(_00988_));
 sky130_fd_sc_hd__nand2_2 _29575_ (.A(_00987_),
    .B(_00988_),
    .Y(_00989_));
 sky130_fd_sc_hd__buf_1 _29576_ (.A(_14352_),
    .X(_00990_));
 sky130_fd_sc_hd__or2_2 _29577_ (.A(_00990_),
    .B(_16922_),
    .X(_00991_));
 sky130_fd_sc_hd__xnor2_2 _29578_ (.A(_00989_),
    .B(_00991_),
    .Y(_00992_));
 sky130_fd_sc_hd__o21a_2 _29579_ (.A1(_00588_),
    .A2(_00590_),
    .B1(_00586_),
    .X(_00993_));
 sky130_fd_sc_hd__xor2_2 _29580_ (.A(_00992_),
    .B(_00993_),
    .X(_00994_));
 sky130_fd_sc_hd__xor2_2 _29581_ (.A(_00984_),
    .B(_00994_),
    .X(_00995_));
 sky130_fd_sc_hd__buf_1 _29582_ (.A(_15835_),
    .X(_00996_));
 sky130_fd_sc_hd__nor2_2 _29583_ (.A(_00996_),
    .B(_00600_),
    .Y(_00998_));
 sky130_fd_sc_hd__buf_1 _29584_ (.A(_13845_),
    .X(_00999_));
 sky130_fd_sc_hd__a22o_2 _29585_ (.A1(_00207_),
    .A2(_00599_),
    .B1(_00998_),
    .B2(_00999_),
    .X(_01000_));
 sky130_fd_sc_hd__o21ba_2 _29586_ (.A1(_00626_),
    .A2(_00628_),
    .B1_N(_00623_),
    .X(_01001_));
 sky130_fd_sc_hd__nor2_2 _29587_ (.A(_15004_),
    .B(_15596_),
    .Y(_01002_));
 sky130_fd_sc_hd__or3b_2 _29588_ (.A(_14988_),
    .B(_16237_),
    .C_N(_01002_),
    .X(_01003_));
 sky130_fd_sc_hd__a2bb2o_2 _29589_ (.A1_N(_14988_),
    .A2_N(_15597_),
    .B1(_15585_),
    .B2(_16292_),
    .X(_01004_));
 sky130_fd_sc_hd__nand2_2 _29590_ (.A(_01003_),
    .B(_01004_),
    .Y(_01005_));
 sky130_fd_sc_hd__nor2_2 _29591_ (.A(_15647_),
    .B(_15835_),
    .Y(_01006_));
 sky130_fd_sc_hd__xnor2_2 _29592_ (.A(_01005_),
    .B(_01006_),
    .Y(_01007_));
 sky130_fd_sc_hd__xnor2_2 _29593_ (.A(_01001_),
    .B(_01007_),
    .Y(_01009_));
 sky130_fd_sc_hd__xnor2_2 _29594_ (.A(_01000_),
    .B(_01009_),
    .Y(_01010_));
 sky130_fd_sc_hd__and2b_2 _29595_ (.A_N(_00598_),
    .B(_00602_),
    .X(_01011_));
 sky130_fd_sc_hd__a21oi_2 _29596_ (.A1(_00596_),
    .A2(_00604_),
    .B1(_01011_),
    .Y(_01012_));
 sky130_fd_sc_hd__or2_2 _29597_ (.A(_01010_),
    .B(_01012_),
    .X(_01013_));
 sky130_fd_sc_hd__nand2_2 _29598_ (.A(_01010_),
    .B(_01012_),
    .Y(_01014_));
 sky130_fd_sc_hd__and3_2 _29599_ (.A(_00995_),
    .B(_01013_),
    .C(_01014_),
    .X(_01015_));
 sky130_fd_sc_hd__and2_2 _29600_ (.A(_01013_),
    .B(_01014_),
    .X(_01016_));
 sky130_fd_sc_hd__nor2_2 _29601_ (.A(_00995_),
    .B(_01016_),
    .Y(_01017_));
 sky130_fd_sc_hd__a211o_2 _29602_ (.A1(_00640_),
    .A2(_00978_),
    .B1(_01015_),
    .C1(_01017_),
    .X(_01018_));
 sky130_fd_sc_hd__o211ai_2 _29603_ (.A1(_01015_),
    .A2(_01017_),
    .B1(_00640_),
    .C1(_00978_),
    .Y(_01020_));
 sky130_fd_sc_hd__o211ai_2 _29604_ (.A1(_00608_),
    .A2(_00611_),
    .B1(_01018_),
    .C1(_01020_),
    .Y(_01021_));
 sky130_fd_sc_hd__a211o_2 _29605_ (.A1(_01018_),
    .A2(_01020_),
    .B1(_00608_),
    .C1(_00611_),
    .X(_01022_));
 sky130_fd_sc_hd__nand3_2 _29606_ (.A(_00643_),
    .B(_00692_),
    .C(_00693_),
    .Y(_01023_));
 sky130_fd_sc_hd__and2b_2 _29607_ (.A_N(_00637_),
    .B(_00635_),
    .X(_01024_));
 sky130_fd_sc_hd__o21ba_2 _29608_ (.A1(_00629_),
    .A2(_00638_),
    .B1_N(_01024_),
    .X(_01025_));
 sky130_fd_sc_hd__nand2_2 _29609_ (.A(_00648_),
    .B(_00654_),
    .Y(_01026_));
 sky130_fd_sc_hd__a21boi_2 _29610_ (.A1(_00646_),
    .A2(_00655_),
    .B1_N(_01026_),
    .Y(_01027_));
 sky130_fd_sc_hd__buf_1 _29611_ (.A(_15169_),
    .X(_01028_));
 sky130_fd_sc_hd__nand2_2 _29612_ (.A(_14410_),
    .B(_00633_),
    .Y(_01029_));
 sky130_fd_sc_hd__o21a_2 _29613_ (.A1(_01028_),
    .A2(_18181_),
    .B1(_01029_),
    .X(_01031_));
 sky130_fd_sc_hd__a31oi_2 _29614_ (.A1(_14606_),
    .A2(_00633_),
    .A3(_00624_),
    .B1(_01031_),
    .Y(_01032_));
 sky130_fd_sc_hd__buf_1 _29615_ (.A(_15617_),
    .X(_01033_));
 sky130_fd_sc_hd__nand2_2 _29616_ (.A(_01033_),
    .B(_15679_),
    .Y(_01034_));
 sky130_fd_sc_hd__xor2_2 _29617_ (.A(_01032_),
    .B(_01034_),
    .X(_01035_));
 sky130_fd_sc_hd__nor2_2 _29618_ (.A(_13893_),
    .B(_16988_),
    .Y(_01036_));
 sky130_fd_sc_hd__nor2_2 _29619_ (.A(_14612_),
    .B(_17007_),
    .Y(_01037_));
 sky130_fd_sc_hd__xnor2_2 _29620_ (.A(_01036_),
    .B(_01037_),
    .Y(_01038_));
 sky130_fd_sc_hd__buf_1 _29621_ (.A(_14391_),
    .X(_01039_));
 sky130_fd_sc_hd__buf_1 _29622_ (.A(_15900_),
    .X(_01040_));
 sky130_fd_sc_hd__nand2_2 _29623_ (.A(_01039_),
    .B(_01040_),
    .Y(_01042_));
 sky130_fd_sc_hd__xnor2_2 _29624_ (.A(_01038_),
    .B(_01042_),
    .Y(_01043_));
 sky130_fd_sc_hd__o21a_2 _29625_ (.A1(_00632_),
    .A2(_00634_),
    .B1(_00630_),
    .X(_01044_));
 sky130_fd_sc_hd__or2_2 _29626_ (.A(_01043_),
    .B(_01044_),
    .X(_01045_));
 sky130_fd_sc_hd__nand2_2 _29627_ (.A(_01043_),
    .B(_01044_),
    .Y(_01046_));
 sky130_fd_sc_hd__nand2_2 _29628_ (.A(_01045_),
    .B(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hd__xor2_2 _29629_ (.A(_01035_),
    .B(_01047_),
    .X(_01048_));
 sky130_fd_sc_hd__xnor2_2 _29630_ (.A(_01027_),
    .B(_01048_),
    .Y(_01049_));
 sky130_fd_sc_hd__xnor2_2 _29631_ (.A(_01025_),
    .B(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__nand3_2 _29632_ (.A(_00656_),
    .B(_00687_),
    .C(_00688_),
    .Y(_01051_));
 sky130_fd_sc_hd__a22o_2 _29633_ (.A1(_00250_),
    .A2(_00650_),
    .B1(_00652_),
    .B2(_17463_),
    .X(_01053_));
 sky130_fd_sc_hd__a21o_2 _29634_ (.A1(_00657_),
    .A2(_00663_),
    .B1(_00660_),
    .X(_01054_));
 sky130_fd_sc_hd__nor2_2 _29635_ (.A(_12852_),
    .B(_17482_),
    .Y(_01055_));
 sky130_fd_sc_hd__and3_2 _29636_ (.A(_14634_),
    .B(_17712_),
    .C(_17713_),
    .X(_01056_));
 sky130_fd_sc_hd__xnor2_2 _29637_ (.A(_01055_),
    .B(_01056_),
    .Y(_01057_));
 sky130_fd_sc_hd__buf_1 _29638_ (.A(_16999_),
    .X(_01058_));
 sky130_fd_sc_hd__or2_2 _29639_ (.A(_14641_),
    .B(_01058_),
    .X(_01059_));
 sky130_fd_sc_hd__xnor2_2 _29640_ (.A(_01057_),
    .B(_01059_),
    .Y(_01060_));
 sky130_fd_sc_hd__xor2_2 _29641_ (.A(_01054_),
    .B(_01060_),
    .X(_01061_));
 sky130_fd_sc_hd__xnor2_2 _29642_ (.A(_01053_),
    .B(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__o22a_2 _29643_ (.A1(_14978_),
    .A2(_00271_),
    .B1(_00666_),
    .B2(_15650_),
    .X(_01064_));
 sky130_fd_sc_hd__a31o_2 _29644_ (.A1(_00661_),
    .A2(_00268_),
    .A3(_00659_),
    .B1(_01064_),
    .X(_01065_));
 sky130_fd_sc_hd__buf_1 _29645_ (.A(_18211_),
    .X(_01066_));
 sky130_fd_sc_hd__nor2_2 _29646_ (.A(_15646_),
    .B(_01066_),
    .Y(_01067_));
 sky130_fd_sc_hd__xnor2_2 _29647_ (.A(_01065_),
    .B(_01067_),
    .Y(_01068_));
 sky130_fd_sc_hd__or2_2 _29648_ (.A(_00278_),
    .B(_00280_),
    .X(_01069_));
 sky130_fd_sc_hd__buf_1 _29649_ (.A(_01069_),
    .X(_01070_));
 sky130_fd_sc_hd__nor2_2 _29650_ (.A(_11794_),
    .B(_01070_),
    .Y(_01071_));
 sky130_fd_sc_hd__or2_2 _29651_ (.A(_00277_),
    .B(_00673_),
    .X(_01072_));
 sky130_fd_sc_hd__or2_2 _29652_ (.A(_18821_),
    .B(_01072_),
    .X(_01073_));
 sky130_fd_sc_hd__a311o_2 _29653_ (.A1(_18446_),
    .A2(_18447_),
    .A3(_18450_),
    .B1(_01073_),
    .C1(_18453_),
    .X(_01075_));
 sky130_fd_sc_hd__nand2_2 _29654_ (.A(_00275_),
    .B(_00672_),
    .Y(_01076_));
 sky130_fd_sc_hd__o2bb2a_2 _29655_ (.A1_N(_00671_),
    .A2_N(_01076_),
    .B1(_01072_),
    .B2(_00279_),
    .X(_01077_));
 sky130_fd_sc_hd__nand2_2 _29656_ (.A(iX[28]),
    .B(iX[60]),
    .Y(_01078_));
 sky130_fd_sc_hd__or2_2 _29657_ (.A(iX[28]),
    .B(iX[60]),
    .X(_01079_));
 sky130_fd_sc_hd__nand2_2 _29658_ (.A(_01078_),
    .B(_01079_),
    .Y(_01080_));
 sky130_fd_sc_hd__a21oi_2 _29659_ (.A1(_01075_),
    .A2(_01077_),
    .B1(_01080_),
    .Y(_01081_));
 sky130_fd_sc_hd__and3_2 _29660_ (.A(_01080_),
    .B(_01075_),
    .C(_01077_),
    .X(_01082_));
 sky130_fd_sc_hd__or3_2 _29661_ (.A(_11576_),
    .B(_01081_),
    .C(_01082_),
    .X(_01083_));
 sky130_fd_sc_hd__or4_4 _29662_ (.A(_11567_),
    .B(_00674_),
    .C(_00675_),
    .D(_01083_),
    .X(_01084_));
 sky130_fd_sc_hd__or2_2 _29663_ (.A(_01081_),
    .B(_01082_),
    .X(_01086_));
 sky130_fd_sc_hd__buf_1 _29664_ (.A(_01086_),
    .X(_01087_));
 sky130_fd_sc_hd__o32ai_2 _29665_ (.A1(_11576_),
    .A2(_00674_),
    .A3(_00675_),
    .B1(_01087_),
    .B2(_11567_),
    .Y(_01088_));
 sky130_fd_sc_hd__nand3_2 _29666_ (.A(_01071_),
    .B(_01084_),
    .C(_01088_),
    .Y(_01089_));
 sky130_fd_sc_hd__a21o_2 _29667_ (.A1(_01084_),
    .A2(_01088_),
    .B1(_01071_),
    .X(_01090_));
 sky130_fd_sc_hd__a21bo_2 _29668_ (.A1(_00667_),
    .A2(_00677_),
    .B1_N(_00676_),
    .X(_01091_));
 sky130_fd_sc_hd__nand3_2 _29669_ (.A(_01089_),
    .B(_01090_),
    .C(_01091_),
    .Y(_01092_));
 sky130_fd_sc_hd__a21o_2 _29670_ (.A1(_01089_),
    .A2(_01090_),
    .B1(_01091_),
    .X(_01093_));
 sky130_fd_sc_hd__nand3_2 _29671_ (.A(_01068_),
    .B(_01092_),
    .C(_01093_),
    .Y(_01094_));
 sky130_fd_sc_hd__a21o_2 _29672_ (.A1(_01092_),
    .A2(_01093_),
    .B1(_01068_),
    .X(_01095_));
 sky130_fd_sc_hd__a21bo_2 _29673_ (.A1(_00665_),
    .A2(_00683_),
    .B1_N(_00682_),
    .X(_01097_));
 sky130_fd_sc_hd__nand3_2 _29674_ (.A(_01094_),
    .B(_01095_),
    .C(_01097_),
    .Y(_01098_));
 sky130_fd_sc_hd__a21o_2 _29675_ (.A1(_01094_),
    .A2(_01095_),
    .B1(_01097_),
    .X(_01099_));
 sky130_fd_sc_hd__and3_2 _29676_ (.A(_01062_),
    .B(_01098_),
    .C(_01099_),
    .X(_01100_));
 sky130_fd_sc_hd__a21oi_2 _29677_ (.A1(_01098_),
    .A2(_01099_),
    .B1(_01062_),
    .Y(_01101_));
 sky130_fd_sc_hd__a211o_2 _29678_ (.A1(_00687_),
    .A2(_01051_),
    .B1(_01100_),
    .C1(_01101_),
    .X(_01102_));
 sky130_fd_sc_hd__o211ai_2 _29679_ (.A1(_01100_),
    .A2(_01101_),
    .B1(_00687_),
    .C1(_01051_),
    .Y(_01103_));
 sky130_fd_sc_hd__and3_4 _29680_ (.A(_01050_),
    .B(_01102_),
    .C(_01103_),
    .X(_01104_));
 sky130_fd_sc_hd__a21oi_2 _29681_ (.A1(_01102_),
    .A2(_01103_),
    .B1(_01050_),
    .Y(_01105_));
 sky130_fd_sc_hd__a211o_2 _29682_ (.A1(_00692_),
    .A2(_01023_),
    .B1(_01104_),
    .C1(_01105_),
    .X(_01106_));
 sky130_fd_sc_hd__o211ai_2 _29683_ (.A1(_01104_),
    .A2(_01105_),
    .B1(_00692_),
    .C1(_01023_),
    .Y(_01108_));
 sky130_fd_sc_hd__nand4_2 _29684_ (.A(_01021_),
    .B(_01022_),
    .C(_01106_),
    .D(_01108_),
    .Y(_01109_));
 sky130_fd_sc_hd__a22o_2 _29685_ (.A1(_01021_),
    .A2(_01022_),
    .B1(_01106_),
    .B2(_01108_),
    .X(_01110_));
 sky130_fd_sc_hd__o211ai_2 _29686_ (.A1(_00696_),
    .A2(_00698_),
    .B1(_01109_),
    .C1(_01110_),
    .Y(_01111_));
 sky130_fd_sc_hd__a211o_2 _29687_ (.A1(_01109_),
    .A2(_01110_),
    .B1(_00696_),
    .C1(_00698_),
    .X(_01112_));
 sky130_fd_sc_hd__and4_4 _29688_ (.A(_00976_),
    .B(_00977_),
    .C(_01111_),
    .D(_01112_),
    .X(_01113_));
 sky130_fd_sc_hd__a22oi_2 _29689_ (.A1(_00976_),
    .A2(_00977_),
    .B1(_01111_),
    .B2(_01112_),
    .Y(_01114_));
 sky130_fd_sc_hd__a211o_2 _29690_ (.A1(_00700_),
    .A2(_00703_),
    .B1(_01113_),
    .C1(_01114_),
    .X(_01115_));
 sky130_fd_sc_hd__o211ai_2 _29691_ (.A1(_01113_),
    .A2(_01114_),
    .B1(_00700_),
    .C1(_00703_),
    .Y(_01116_));
 sky130_fd_sc_hd__o211ai_2 _29692_ (.A1(_00571_),
    .A2(_00574_),
    .B1(_01115_),
    .C1(_01116_),
    .Y(_01117_));
 sky130_fd_sc_hd__a211o_2 _29693_ (.A1(_01115_),
    .A2(_01116_),
    .B1(_00571_),
    .C1(_00574_),
    .X(_01119_));
 sky130_fd_sc_hd__o211ai_2 _29694_ (.A1(_00705_),
    .A2(_00928_),
    .B1(_01117_),
    .C1(_01119_),
    .Y(_01120_));
 sky130_fd_sc_hd__a211o_2 _29695_ (.A1(_01117_),
    .A2(_01119_),
    .B1(_00705_),
    .C1(_00928_),
    .X(_01121_));
 sky130_fd_sc_hd__nand2_2 _29696_ (.A(_01120_),
    .B(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__xnor2_2 _29697_ (.A(_00709_),
    .B(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__or4_4 _29698_ (.A(_18497_),
    .B(_18498_),
    .C(_18849_),
    .D(_18850_),
    .X(_01124_));
 sky130_fd_sc_hd__or4_4 _29699_ (.A(_00314_),
    .B(_00711_),
    .C(_00712_),
    .D(_01124_),
    .X(_01125_));
 sky130_fd_sc_hd__a21o_2 _29700_ (.A1(_18315_),
    .A2(_18318_),
    .B1(_01125_),
    .X(_01126_));
 sky130_fd_sc_hd__or2_2 _29701_ (.A(_18849_),
    .B(_00315_),
    .X(_01127_));
 sky130_fd_sc_hd__nand2_2 _29702_ (.A(_00709_),
    .B(_00710_),
    .Y(_01128_));
 sky130_fd_sc_hd__o21ba_2 _29703_ (.A1(_00523_),
    .A2(_01128_),
    .B1_N(_00711_),
    .X(_01130_));
 sky130_fd_sc_hd__o31a_2 _29704_ (.A1(_00314_),
    .A2(_00714_),
    .A3(_01127_),
    .B1(_01130_),
    .X(_01131_));
 sky130_fd_sc_hd__and2_2 _29705_ (.A(_01126_),
    .B(_01131_),
    .X(_01132_));
 sky130_fd_sc_hd__xnor2_2 _29706_ (.A(_01123_),
    .B(_01132_),
    .Y(_01133_));
 sky130_fd_sc_hd__a211o_2 _29707_ (.A1(_00466_),
    .A2(_00467_),
    .B1(_00880_),
    .C1(_00874_),
    .X(_01134_));
 sky130_fd_sc_hd__o21ba_2 _29708_ (.A1(_00875_),
    .A2(_00873_),
    .B1_N(_00877_),
    .X(_01135_));
 sky130_fd_sc_hd__inv_2 _29709_ (.A(_00860_),
    .Y(_01136_));
 sky130_fd_sc_hd__nand2_2 _29710_ (.A(_00785_),
    .B(_00786_),
    .Y(_01137_));
 sky130_fd_sc_hd__and3_2 _29711_ (.A(_00751_),
    .B(_00752_),
    .C(_00754_),
    .X(_01138_));
 sky130_fd_sc_hd__or2b_2 _29712_ (.A(_00728_),
    .B_N(_00727_),
    .X(_01139_));
 sky130_fd_sc_hd__nand2_2 _29713_ (.A(_00729_),
    .B(_00737_),
    .Y(_01141_));
 sky130_fd_sc_hd__and4_2 _29714_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[57]),
    .D(iX[58]),
    .X(_01142_));
 sky130_fd_sc_hd__a22oi_2 _29715_ (.A1(iY[35]),
    .A2(iX[57]),
    .B1(iX[58]),
    .B2(iY[34]),
    .Y(_01143_));
 sky130_fd_sc_hd__nor2_2 _29716_ (.A(_01142_),
    .B(_01143_),
    .Y(_01144_));
 sky130_fd_sc_hd__nand2_2 _29717_ (.A(iY[33]),
    .B(iX[59]),
    .Y(_01145_));
 sky130_fd_sc_hd__xnor2_2 _29718_ (.A(_01144_),
    .B(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hd__o21ba_2 _29719_ (.A1(_00723_),
    .A2(_00726_),
    .B1_N(_00722_),
    .X(_01147_));
 sky130_fd_sc_hd__xnor2_2 _29720_ (.A(_01146_),
    .B(_01147_),
    .Y(_01148_));
 sky130_fd_sc_hd__and4_2 _29721_ (.A(iY[32]),
    .B(iY[36]),
    .C(iX[56]),
    .D(iX[60]),
    .X(_01149_));
 sky130_fd_sc_hd__a22oi_2 _29722_ (.A1(iY[36]),
    .A2(iX[56]),
    .B1(iX[60]),
    .B2(iY[32]),
    .Y(_01150_));
 sky130_fd_sc_hd__o2bb2a_2 _29723_ (.A1_N(iY[37]),
    .A2_N(iX[55]),
    .B1(_01149_),
    .B2(_01150_),
    .X(_01152_));
 sky130_fd_sc_hd__and4bb_2 _29724_ (.A_N(_01149_),
    .B_N(_01150_),
    .C(iY[37]),
    .D(iX[55]),
    .X(_01153_));
 sky130_fd_sc_hd__nor2_2 _29725_ (.A(_01152_),
    .B(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__xnor2_2 _29726_ (.A(_01148_),
    .B(_01154_),
    .Y(_01155_));
 sky130_fd_sc_hd__a21o_2 _29727_ (.A1(_01139_),
    .A2(_01141_),
    .B1(_01155_),
    .X(_01156_));
 sky130_fd_sc_hd__nand3_2 _29728_ (.A(_01139_),
    .B(_01141_),
    .C(_01155_),
    .Y(_01157_));
 sky130_fd_sc_hd__o21ba_2 _29729_ (.A1(_00744_),
    .A2(_00747_),
    .B1_N(_00743_),
    .X(_01158_));
 sky130_fd_sc_hd__and3_2 _29730_ (.A(iY[32]),
    .B(iX[55]),
    .C(_00730_),
    .X(_01159_));
 sky130_fd_sc_hd__and4_2 _29731_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[53]),
    .D(iX[54]),
    .X(_01160_));
 sky130_fd_sc_hd__a22oi_2 _29732_ (.A1(iY[39]),
    .A2(iX[53]),
    .B1(iX[54]),
    .B2(iY[38]),
    .Y(_01161_));
 sky130_fd_sc_hd__nor2_2 _29733_ (.A(_01160_),
    .B(_01161_),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2_2 _29734_ (.A(iY[40]),
    .B(iX[52]),
    .Y(_01164_));
 sky130_fd_sc_hd__xnor2_2 _29735_ (.A(_01163_),
    .B(_01164_),
    .Y(_01165_));
 sky130_fd_sc_hd__o21ai_2 _29736_ (.A1(_01159_),
    .A2(_00736_),
    .B1(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__or3_2 _29737_ (.A(_01159_),
    .B(_00736_),
    .C(_01165_),
    .X(_01167_));
 sky130_fd_sc_hd__and2_2 _29738_ (.A(_01166_),
    .B(_01167_),
    .X(_01168_));
 sky130_fd_sc_hd__xnor2_2 _29739_ (.A(_01158_),
    .B(_01168_),
    .Y(_01169_));
 sky130_fd_sc_hd__nand3_2 _29740_ (.A(_01156_),
    .B(_01157_),
    .C(_01169_),
    .Y(_01170_));
 sky130_fd_sc_hd__a21o_2 _29741_ (.A1(_01156_),
    .A2(_01157_),
    .B1(_01169_),
    .X(_01171_));
 sky130_fd_sc_hd__nand2_2 _29742_ (.A(_01170_),
    .B(_01171_),
    .Y(_01172_));
 sky130_fd_sc_hd__nand2_2 _29743_ (.A(_00739_),
    .B(_00751_),
    .Y(_01174_));
 sky130_fd_sc_hd__xnor2_2 _29744_ (.A(_01172_),
    .B(_01174_),
    .Y(_01175_));
 sky130_fd_sc_hd__and2b_2 _29745_ (.A_N(_00771_),
    .B(_00770_),
    .X(_01176_));
 sky130_fd_sc_hd__or2b_2 _29746_ (.A(_00742_),
    .B_N(_00748_),
    .X(_01177_));
 sky130_fd_sc_hd__or2b_2 _29747_ (.A(_00741_),
    .B_N(_00749_),
    .X(_01178_));
 sky130_fd_sc_hd__and4_2 _29748_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[47]),
    .D(iX[48]),
    .X(_01179_));
 sky130_fd_sc_hd__a22oi_2 _29749_ (.A1(iY[45]),
    .A2(iX[47]),
    .B1(iX[48]),
    .B2(iY[44]),
    .Y(_01180_));
 sky130_fd_sc_hd__nor2_2 _29750_ (.A(_01179_),
    .B(_01180_),
    .Y(_01181_));
 sky130_fd_sc_hd__nand2_2 _29751_ (.A(iX[46]),
    .B(iY[46]),
    .Y(_01182_));
 sky130_fd_sc_hd__xnor2_2 _29752_ (.A(_01181_),
    .B(_01182_),
    .Y(_01183_));
 sky130_fd_sc_hd__and4_2 _29753_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[50]),
    .D(iX[51]),
    .X(_01185_));
 sky130_fd_sc_hd__a22oi_2 _29754_ (.A1(iY[42]),
    .A2(iX[50]),
    .B1(iX[51]),
    .B2(iY[41]),
    .Y(_01186_));
 sky130_fd_sc_hd__nor2_2 _29755_ (.A(_01185_),
    .B(_01186_),
    .Y(_01187_));
 sky130_fd_sc_hd__nand2_2 _29756_ (.A(iY[43]),
    .B(iX[49]),
    .Y(_01188_));
 sky130_fd_sc_hd__xnor2_2 _29757_ (.A(_01187_),
    .B(_01188_),
    .Y(_01189_));
 sky130_fd_sc_hd__o21ba_2 _29758_ (.A1(_00766_),
    .A2(_00769_),
    .B1_N(_00765_),
    .X(_01190_));
 sky130_fd_sc_hd__xnor2_2 _29759_ (.A(_01189_),
    .B(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__and2_2 _29760_ (.A(_01183_),
    .B(_01191_),
    .X(_01192_));
 sky130_fd_sc_hd__nor2_2 _29761_ (.A(_01183_),
    .B(_01191_),
    .Y(_01193_));
 sky130_fd_sc_hd__or2_2 _29762_ (.A(_01192_),
    .B(_01193_),
    .X(_01194_));
 sky130_fd_sc_hd__a21o_2 _29763_ (.A1(_01177_),
    .A2(_01178_),
    .B1(_01194_),
    .X(_01196_));
 sky130_fd_sc_hd__nand3_2 _29764_ (.A(_01177_),
    .B(_01178_),
    .C(_01194_),
    .Y(_01197_));
 sky130_fd_sc_hd__o211ai_2 _29765_ (.A1(_01176_),
    .A2(_00773_),
    .B1(_01196_),
    .C1(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hd__a211o_2 _29766_ (.A1(_01196_),
    .A2(_01197_),
    .B1(_01176_),
    .C1(_00773_),
    .X(_01199_));
 sky130_fd_sc_hd__and3_2 _29767_ (.A(_01175_),
    .B(_01198_),
    .C(_01199_),
    .X(_01200_));
 sky130_fd_sc_hd__inv_2 _29768_ (.A(_01200_),
    .Y(_01201_));
 sky130_fd_sc_hd__a21o_2 _29769_ (.A1(_01198_),
    .A2(_01199_),
    .B1(_01175_),
    .X(_01202_));
 sky130_fd_sc_hd__o211ai_2 _29770_ (.A1(_01138_),
    .A2(_00783_),
    .B1(_01201_),
    .C1(_01202_),
    .Y(_01203_));
 sky130_fd_sc_hd__a211o_2 _29771_ (.A1(_01201_),
    .A2(_01202_),
    .B1(_01138_),
    .C1(_00783_),
    .X(_01204_));
 sky130_fd_sc_hd__nand2_2 _29772_ (.A(_01203_),
    .B(_01204_),
    .Y(_01205_));
 sky130_fd_sc_hd__a21o_2 _29773_ (.A1(_00805_),
    .A2(_00413_),
    .B1(_00816_),
    .X(_01207_));
 sky130_fd_sc_hd__and4_2 _29774_ (.A(iX[38]),
    .B(iX[39]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_01208_));
 sky130_fd_sc_hd__a22oi_2 _29775_ (.A1(iX[39]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[38]),
    .Y(_01209_));
 sky130_fd_sc_hd__nor2_2 _29776_ (.A(_01208_),
    .B(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__nand2_2 _29777_ (.A(iX[37]),
    .B(iY[55]),
    .Y(_01211_));
 sky130_fd_sc_hd__xnor2_2 _29778_ (.A(_01210_),
    .B(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hd__and4_2 _29779_ (.A(iX[41]),
    .B(iX[42]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_01213_));
 sky130_fd_sc_hd__a22oi_2 _29780_ (.A1(iX[42]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[41]),
    .Y(_01214_));
 sky130_fd_sc_hd__nor2_2 _29781_ (.A(_01213_),
    .B(_01214_),
    .Y(_01215_));
 sky130_fd_sc_hd__nand2_2 _29782_ (.A(iX[40]),
    .B(iY[52]),
    .Y(_01216_));
 sky130_fd_sc_hd__xnor2_2 _29783_ (.A(_01215_),
    .B(_01216_),
    .Y(_01218_));
 sky130_fd_sc_hd__o21ba_2 _29784_ (.A1(_00795_),
    .A2(_00797_),
    .B1_N(_00794_),
    .X(_01219_));
 sky130_fd_sc_hd__xnor2_2 _29785_ (.A(_01218_),
    .B(_01219_),
    .Y(_01220_));
 sky130_fd_sc_hd__and2_2 _29786_ (.A(_01212_),
    .B(_01220_),
    .X(_01221_));
 sky130_fd_sc_hd__nor2_2 _29787_ (.A(_01212_),
    .B(_01220_),
    .Y(_01222_));
 sky130_fd_sc_hd__or2_2 _29788_ (.A(_01221_),
    .B(_01222_),
    .X(_01223_));
 sky130_fd_sc_hd__or3_2 _29789_ (.A(_00806_),
    .B(_00809_),
    .C(_00810_),
    .X(_01224_));
 sky130_fd_sc_hd__o21ba_2 _29790_ (.A1(_00761_),
    .A2(_00763_),
    .B1_N(_00760_),
    .X(_01225_));
 sky130_fd_sc_hd__and4_2 _29791_ (.A(iX[44]),
    .B(iX[45]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_01226_));
 sky130_fd_sc_hd__a22oi_2 _29792_ (.A1(iX[45]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[44]),
    .Y(_01227_));
 sky130_fd_sc_hd__nand2_2 _29793_ (.A(iX[43]),
    .B(iY[49]),
    .Y(_01229_));
 sky130_fd_sc_hd__o21a_2 _29794_ (.A1(_01226_),
    .A2(_01227_),
    .B1(_01229_),
    .X(_01230_));
 sky130_fd_sc_hd__nor3_2 _29795_ (.A(_01226_),
    .B(_01227_),
    .C(_01229_),
    .Y(_01231_));
 sky130_fd_sc_hd__nor2_2 _29796_ (.A(_01230_),
    .B(_01231_),
    .Y(_01232_));
 sky130_fd_sc_hd__xnor2_2 _29797_ (.A(_01225_),
    .B(_01232_),
    .Y(_01233_));
 sky130_fd_sc_hd__o21ai_2 _29798_ (.A1(_00807_),
    .A2(_00809_),
    .B1(_01233_),
    .Y(_01234_));
 sky130_fd_sc_hd__or3_2 _29799_ (.A(_00807_),
    .B(_00809_),
    .C(_01233_),
    .X(_01235_));
 sky130_fd_sc_hd__nand2_2 _29800_ (.A(_01234_),
    .B(_01235_),
    .Y(_01236_));
 sky130_fd_sc_hd__a21oi_2 _29801_ (.A1(_01224_),
    .A2(_00814_),
    .B1(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__and3_2 _29802_ (.A(_01224_),
    .B(_00814_),
    .C(_01236_),
    .X(_01238_));
 sky130_fd_sc_hd__or3_2 _29803_ (.A(_01223_),
    .B(_01237_),
    .C(_01238_),
    .X(_01240_));
 sky130_fd_sc_hd__o21ai_2 _29804_ (.A1(_01237_),
    .A2(_01238_),
    .B1(_01223_),
    .Y(_01241_));
 sky130_fd_sc_hd__nand2_2 _29805_ (.A(_01240_),
    .B(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hd__a21oi_2 _29806_ (.A1(_00776_),
    .A2(_00780_),
    .B1(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__and3_2 _29807_ (.A(_00776_),
    .B(_00780_),
    .C(_01242_),
    .X(_01244_));
 sky130_fd_sc_hd__a211oi_2 _29808_ (.A1(_01207_),
    .A2(_00819_),
    .B1(_01243_),
    .C1(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__o211a_2 _29809_ (.A1(_01243_),
    .A2(_01244_),
    .B1(_01207_),
    .C1(_00819_),
    .X(_01246_));
 sky130_fd_sc_hd__or3_2 _29810_ (.A(_01205_),
    .B(_01245_),
    .C(_01246_),
    .X(_01247_));
 sky130_fd_sc_hd__inv_2 _29811_ (.A(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hd__o21a_2 _29812_ (.A1(_01245_),
    .A2(_01246_),
    .B1(_01205_),
    .X(_01249_));
 sky130_fd_sc_hd__a211o_2 _29813_ (.A1(_01137_),
    .A2(_00827_),
    .B1(_01248_),
    .C1(_01249_),
    .X(_01251_));
 sky130_fd_sc_hd__inv_2 _29814_ (.A(_01251_),
    .Y(_01252_));
 sky130_fd_sc_hd__o211a_2 _29815_ (.A1(_01248_),
    .A2(_01249_),
    .B1(_01137_),
    .C1(_00827_),
    .X(_01253_));
 sky130_fd_sc_hd__nor2_2 _29816_ (.A(_01252_),
    .B(_01253_),
    .Y(_01254_));
 sky130_fd_sc_hd__a22o_2 _29817_ (.A1(iX[33]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[32]),
    .X(_01255_));
 sky130_fd_sc_hd__and4_2 _29818_ (.A(iX[33]),
    .B(iX[32]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_01256_));
 sky130_fd_sc_hd__inv_2 _29819_ (.A(_01256_),
    .Y(_01257_));
 sky130_fd_sc_hd__or2b_2 _29820_ (.A(_00835_),
    .B_N(_00840_),
    .X(_01258_));
 sky130_fd_sc_hd__or2b_2 _29821_ (.A(_00833_),
    .B_N(_00841_),
    .X(_01259_));
 sky130_fd_sc_hd__and2b_2 _29822_ (.A_N(_00799_),
    .B(_00798_),
    .X(_01260_));
 sky130_fd_sc_hd__o21ba_2 _29823_ (.A1(_00837_),
    .A2(_00839_),
    .B1_N(_00836_),
    .X(_01262_));
 sky130_fd_sc_hd__o21ba_2 _29824_ (.A1(_00789_),
    .A2(_00792_),
    .B1_N(_00788_),
    .X(_01263_));
 sky130_fd_sc_hd__and4_2 _29825_ (.A(iX[35]),
    .B(iX[36]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_01264_));
 sky130_fd_sc_hd__a22oi_2 _29826_ (.A1(iX[36]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[35]),
    .Y(_01265_));
 sky130_fd_sc_hd__nor2_2 _29827_ (.A(_01264_),
    .B(_01265_),
    .Y(_01266_));
 sky130_fd_sc_hd__nand2_2 _29828_ (.A(iX[34]),
    .B(iY[58]),
    .Y(_01267_));
 sky130_fd_sc_hd__xnor2_2 _29829_ (.A(_01266_),
    .B(_01267_),
    .Y(_01268_));
 sky130_fd_sc_hd__xnor2_2 _29830_ (.A(_01263_),
    .B(_01268_),
    .Y(_01269_));
 sky130_fd_sc_hd__xnor2_2 _29831_ (.A(_01262_),
    .B(_01269_),
    .Y(_01270_));
 sky130_fd_sc_hd__o21a_2 _29832_ (.A1(_01260_),
    .A2(_00802_),
    .B1(_01270_),
    .X(_01271_));
 sky130_fd_sc_hd__nor3_2 _29833_ (.A(_01260_),
    .B(_00802_),
    .C(_01270_),
    .Y(_01273_));
 sky130_fd_sc_hd__a211oi_2 _29834_ (.A1(_01258_),
    .A2(_01259_),
    .B1(_01271_),
    .C1(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hd__o211a_2 _29835_ (.A1(_01271_),
    .A2(_01273_),
    .B1(_01258_),
    .C1(_01259_),
    .X(_01275_));
 sky130_fd_sc_hd__nor2_2 _29836_ (.A(_00843_),
    .B(_00848_),
    .Y(_01276_));
 sky130_fd_sc_hd__or3_2 _29837_ (.A(_01274_),
    .B(_01275_),
    .C(_01276_),
    .X(_01277_));
 sky130_fd_sc_hd__o21ai_2 _29838_ (.A1(_01274_),
    .A2(_01275_),
    .B1(_01276_),
    .Y(_01278_));
 sky130_fd_sc_hd__nand4_2 _29839_ (.A(_01255_),
    .B(_01257_),
    .C(_01277_),
    .D(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hd__a22o_2 _29840_ (.A1(_01255_),
    .A2(_01257_),
    .B1(_01277_),
    .B2(_01278_),
    .X(_01280_));
 sky130_fd_sc_hd__o211a_2 _29841_ (.A1(_00821_),
    .A2(_00825_),
    .B1(_01279_),
    .C1(_01280_),
    .X(_01281_));
 sky130_fd_sc_hd__a211oi_2 _29842_ (.A1(_01279_),
    .A2(_01280_),
    .B1(_00821_),
    .C1(_00825_),
    .Y(_01282_));
 sky130_fd_sc_hd__a211oi_2 _29843_ (.A1(_00852_),
    .A2(_00857_),
    .B1(_01281_),
    .C1(_01282_),
    .Y(_01284_));
 sky130_fd_sc_hd__o211a_2 _29844_ (.A1(_01281_),
    .A2(_01282_),
    .B1(_00852_),
    .C1(_00857_),
    .X(_01285_));
 sky130_fd_sc_hd__nor2_2 _29845_ (.A(_01284_),
    .B(_01285_),
    .Y(_01286_));
 sky130_fd_sc_hd__xnor2_2 _29846_ (.A(_01254_),
    .B(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__a21oi_2 _29847_ (.A1(_00830_),
    .A2(_00864_),
    .B1(_01287_),
    .Y(_01288_));
 sky130_fd_sc_hd__and3_2 _29848_ (.A(_00830_),
    .B(_00864_),
    .C(_01287_),
    .X(_01289_));
 sky130_fd_sc_hd__a211oi_2 _29849_ (.A1(_01136_),
    .A2(_00863_),
    .B1(_01288_),
    .C1(_01289_),
    .Y(_01290_));
 sky130_fd_sc_hd__o211a_2 _29850_ (.A1(_01288_),
    .A2(_01289_),
    .B1(_01136_),
    .C1(_00863_),
    .X(_01291_));
 sky130_fd_sc_hd__or2_2 _29851_ (.A(_01290_),
    .B(_01291_),
    .X(_01292_));
 sky130_fd_sc_hd__nand2_2 _29852_ (.A(_00866_),
    .B(_00869_),
    .Y(_01293_));
 sky130_fd_sc_hd__xnor2_2 _29853_ (.A(_01292_),
    .B(_01293_),
    .Y(_01295_));
 sky130_fd_sc_hd__xor2_2 _29854_ (.A(_00871_),
    .B(_01295_),
    .X(_01296_));
 sky130_fd_sc_hd__a21oi_2 _29855_ (.A1(_01134_),
    .A2(_01135_),
    .B1(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__and3_2 _29856_ (.A(_01134_),
    .B(_01296_),
    .C(_01135_),
    .X(_01298_));
 sky130_fd_sc_hd__nor2_2 _29857_ (.A(_01297_),
    .B(_01298_),
    .Y(_01299_));
 sky130_fd_sc_hd__xor2_2 _29858_ (.A(_01133_),
    .B(_01299_),
    .X(_01300_));
 sky130_fd_sc_hd__nand2_2 _29859_ (.A(_10671_),
    .B(_01300_),
    .Y(_01301_));
 sky130_fd_sc_hd__or2_2 _29860_ (.A(_10671_),
    .B(_01300_),
    .X(_01302_));
 sky130_fd_sc_hd__nand2_2 _29861_ (.A(_01301_),
    .B(_01302_),
    .Y(_01303_));
 sky130_fd_sc_hd__and2b_2 _29862_ (.A_N(_00884_),
    .B(_00885_),
    .X(_01304_));
 sky130_fd_sc_hd__xnor2_2 _29863_ (.A(_01303_),
    .B(_01304_),
    .Y(_01306_));
 sky130_fd_sc_hd__xnor2_2 _29864_ (.A(_00927_),
    .B(_01306_),
    .Y(_01307_));
 sky130_fd_sc_hd__nand2_2 _29865_ (.A(_00924_),
    .B(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__or2_2 _29866_ (.A(_00924_),
    .B(_01307_),
    .X(_01309_));
 sky130_fd_sc_hd__nand2_2 _29867_ (.A(_01308_),
    .B(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__a21bo_2 _29868_ (.A1(_00522_),
    .A2(_00895_),
    .B1_N(_00482_),
    .X(_01311_));
 sky130_fd_sc_hd__o21ai_2 _29869_ (.A1(_00522_),
    .A2(_00895_),
    .B1(_01311_),
    .Y(_01312_));
 sky130_fd_sc_hd__or2_2 _29870_ (.A(_00100_),
    .B(_01312_),
    .X(_01313_));
 sky130_fd_sc_hd__and2_2 _29871_ (.A(_00485_),
    .B(_00896_),
    .X(_01314_));
 sky130_fd_sc_hd__o22a_2 _29872_ (.A1(_00097_),
    .A2(_01313_),
    .B1(_01314_),
    .B2(_01312_),
    .X(_01315_));
 sky130_fd_sc_hd__xnor2_2 _29873_ (.A(_01310_),
    .B(_01315_),
    .Y(oO[60]));
 sky130_fd_sc_hd__and2b_2 _29874_ (.A_N(_00917_),
    .B(_00916_),
    .X(_01317_));
 sky130_fd_sc_hd__a21oi_2 _29875_ (.A1(_00103_),
    .A2(_00902_),
    .B1(_00491_),
    .Y(_01318_));
 sky130_fd_sc_hd__and3_2 _29876_ (.A(iY[30]),
    .B(iX[31]),
    .C(_01318_),
    .X(_01319_));
 sky130_fd_sc_hd__a21oi_2 _29877_ (.A1(iY[30]),
    .A2(iX[31]),
    .B1(_01318_),
    .Y(_01320_));
 sky130_fd_sc_hd__or2_2 _29878_ (.A(_01319_),
    .B(_01320_),
    .X(_01321_));
 sky130_fd_sc_hd__nand2_2 _29879_ (.A(iX[30]),
    .B(iY[31]),
    .Y(_01322_));
 sky130_fd_sc_hd__xor2_2 _29880_ (.A(_01321_),
    .B(_01322_),
    .X(_01323_));
 sky130_fd_sc_hd__xnor2_2 _29881_ (.A(_00911_),
    .B(_01323_),
    .Y(_01324_));
 sky130_fd_sc_hd__o21ba_2 _29882_ (.A1(_00903_),
    .A2(_00904_),
    .B1_N(_00908_),
    .X(_01325_));
 sky130_fd_sc_hd__xnor2_2 _29883_ (.A(_01324_),
    .B(_01325_),
    .Y(_01327_));
 sky130_fd_sc_hd__o21ai_2 _29884_ (.A1(_00914_),
    .A2(_01317_),
    .B1(_01327_),
    .Y(_01328_));
 sky130_fd_sc_hd__or3_2 _29885_ (.A(_00914_),
    .B(_01317_),
    .C(_01327_),
    .X(_01329_));
 sky130_fd_sc_hd__and2_2 _29886_ (.A(_01328_),
    .B(_01329_),
    .X(_01330_));
 sky130_fd_sc_hd__inv_2 _29887_ (.A(_01330_),
    .Y(_01331_));
 sky130_fd_sc_hd__inv_2 _29888_ (.A(_00921_),
    .Y(_01332_));
 sky130_fd_sc_hd__a21oi_2 _29889_ (.A1(_01332_),
    .A2(_00923_),
    .B1(_00919_),
    .Y(_01333_));
 sky130_fd_sc_hd__xnor2_2 _29890_ (.A(_01331_),
    .B(_01333_),
    .Y(_01334_));
 sky130_fd_sc_hd__inv_2 _29891_ (.A(_01334_),
    .Y(_01335_));
 sky130_fd_sc_hd__or2_2 _29892_ (.A(_01133_),
    .B(_01299_),
    .X(_01336_));
 sky130_fd_sc_hd__and2b_2 _29893_ (.A_N(_01292_),
    .B(_01293_),
    .X(_01338_));
 sky130_fd_sc_hd__and3_2 _29894_ (.A(_01170_),
    .B(_01171_),
    .C(_01174_),
    .X(_01339_));
 sky130_fd_sc_hd__and2b_2 _29895_ (.A_N(_01190_),
    .B(_01189_),
    .X(_01340_));
 sky130_fd_sc_hd__or2b_2 _29896_ (.A(_01158_),
    .B_N(_01168_),
    .X(_01341_));
 sky130_fd_sc_hd__and4_2 _29897_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[48]),
    .D(iX[49]),
    .X(_01342_));
 sky130_fd_sc_hd__a22oi_2 _29898_ (.A1(iY[45]),
    .A2(iX[48]),
    .B1(iX[49]),
    .B2(iY[44]),
    .Y(_01343_));
 sky130_fd_sc_hd__nor2_2 _29899_ (.A(_01342_),
    .B(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__nand2_2 _29900_ (.A(iY[46]),
    .B(iX[47]),
    .Y(_01345_));
 sky130_fd_sc_hd__xnor2_2 _29901_ (.A(_01344_),
    .B(_01345_),
    .Y(_01346_));
 sky130_fd_sc_hd__and4_2 _29902_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[51]),
    .D(iX[52]),
    .X(_01347_));
 sky130_fd_sc_hd__a22oi_2 _29903_ (.A1(iY[42]),
    .A2(iX[51]),
    .B1(iX[52]),
    .B2(iY[41]),
    .Y(_01349_));
 sky130_fd_sc_hd__nor2_2 _29904_ (.A(_01347_),
    .B(_01349_),
    .Y(_01350_));
 sky130_fd_sc_hd__nand2_2 _29905_ (.A(iY[43]),
    .B(iX[50]),
    .Y(_01351_));
 sky130_fd_sc_hd__xnor2_2 _29906_ (.A(_01350_),
    .B(_01351_),
    .Y(_01352_));
 sky130_fd_sc_hd__o21ba_2 _29907_ (.A1(_01186_),
    .A2(_01188_),
    .B1_N(_01185_),
    .X(_01353_));
 sky130_fd_sc_hd__xnor2_2 _29908_ (.A(_01352_),
    .B(_01353_),
    .Y(_01354_));
 sky130_fd_sc_hd__and2_2 _29909_ (.A(_01346_),
    .B(_01354_),
    .X(_01355_));
 sky130_fd_sc_hd__nor2_2 _29910_ (.A(_01346_),
    .B(_01354_),
    .Y(_01356_));
 sky130_fd_sc_hd__or2_2 _29911_ (.A(_01355_),
    .B(_01356_),
    .X(_01357_));
 sky130_fd_sc_hd__a21o_2 _29912_ (.A1(_01166_),
    .A2(_01341_),
    .B1(_01357_),
    .X(_01358_));
 sky130_fd_sc_hd__nand3_2 _29913_ (.A(_01166_),
    .B(_01341_),
    .C(_01357_),
    .Y(_01360_));
 sky130_fd_sc_hd__o211ai_2 _29914_ (.A1(_01340_),
    .A2(_01192_),
    .B1(_01358_),
    .C1(_01360_),
    .Y(_01361_));
 sky130_fd_sc_hd__a211o_2 _29915_ (.A1(_01358_),
    .A2(_01360_),
    .B1(_01340_),
    .C1(_01192_),
    .X(_01362_));
 sky130_fd_sc_hd__or2b_2 _29916_ (.A(_01147_),
    .B_N(_01146_),
    .X(_01363_));
 sky130_fd_sc_hd__nand2_2 _29917_ (.A(_01148_),
    .B(_01154_),
    .Y(_01364_));
 sky130_fd_sc_hd__and4_2 _29918_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[58]),
    .D(iX[59]),
    .X(_01365_));
 sky130_fd_sc_hd__a22oi_2 _29919_ (.A1(iY[35]),
    .A2(iX[58]),
    .B1(iX[59]),
    .B2(iY[34]),
    .Y(_01366_));
 sky130_fd_sc_hd__nor2_2 _29920_ (.A(_01365_),
    .B(_01366_),
    .Y(_01367_));
 sky130_fd_sc_hd__nand2_2 _29921_ (.A(iY[33]),
    .B(iX[60]),
    .Y(_01368_));
 sky130_fd_sc_hd__xnor2_2 _29922_ (.A(_01367_),
    .B(_01368_),
    .Y(_01369_));
 sky130_fd_sc_hd__o21ba_2 _29923_ (.A1(_01143_),
    .A2(_01145_),
    .B1_N(_01142_),
    .X(_01371_));
 sky130_fd_sc_hd__xnor2_2 _29924_ (.A(_01369_),
    .B(_01371_),
    .Y(_01372_));
 sky130_fd_sc_hd__and2_2 _29925_ (.A(iY[36]),
    .B(iX[61]),
    .X(_01373_));
 sky130_fd_sc_hd__and3_2 _29926_ (.A(iY[32]),
    .B(iX[57]),
    .C(_01373_),
    .X(_01374_));
 sky130_fd_sc_hd__a22oi_2 _29927_ (.A1(iY[36]),
    .A2(iX[57]),
    .B1(iX[61]),
    .B2(iY[32]),
    .Y(_01375_));
 sky130_fd_sc_hd__o2bb2a_2 _29928_ (.A1_N(iY[37]),
    .A2_N(iX[56]),
    .B1(_01374_),
    .B2(_01375_),
    .X(_01376_));
 sky130_fd_sc_hd__and4bb_2 _29929_ (.A_N(_01374_),
    .B_N(_01375_),
    .C(iY[37]),
    .D(iX[56]),
    .X(_01377_));
 sky130_fd_sc_hd__nor2_2 _29930_ (.A(_01376_),
    .B(_01377_),
    .Y(_01378_));
 sky130_fd_sc_hd__xnor2_2 _29931_ (.A(_01372_),
    .B(_01378_),
    .Y(_01379_));
 sky130_fd_sc_hd__a21o_2 _29932_ (.A1(_01363_),
    .A2(_01364_),
    .B1(_01379_),
    .X(_01380_));
 sky130_fd_sc_hd__nand3_2 _29933_ (.A(_01363_),
    .B(_01364_),
    .C(_01379_),
    .Y(_01382_));
 sky130_fd_sc_hd__o21ba_2 _29934_ (.A1(_01161_),
    .A2(_01164_),
    .B1_N(_01160_),
    .X(_01383_));
 sky130_fd_sc_hd__and4_2 _29935_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[54]),
    .D(iX[55]),
    .X(_01384_));
 sky130_fd_sc_hd__a22oi_2 _29936_ (.A1(iY[39]),
    .A2(iX[54]),
    .B1(iX[55]),
    .B2(iY[38]),
    .Y(_01385_));
 sky130_fd_sc_hd__nor2_2 _29937_ (.A(_01384_),
    .B(_01385_),
    .Y(_01386_));
 sky130_fd_sc_hd__nand2_2 _29938_ (.A(iY[40]),
    .B(iX[53]),
    .Y(_01387_));
 sky130_fd_sc_hd__xnor2_2 _29939_ (.A(_01386_),
    .B(_01387_),
    .Y(_01388_));
 sky130_fd_sc_hd__o21ai_2 _29940_ (.A1(_01149_),
    .A2(_01153_),
    .B1(_01388_),
    .Y(_01389_));
 sky130_fd_sc_hd__or3_2 _29941_ (.A(_01149_),
    .B(_01153_),
    .C(_01388_),
    .X(_01390_));
 sky130_fd_sc_hd__and2_2 _29942_ (.A(_01389_),
    .B(_01390_),
    .X(_01391_));
 sky130_fd_sc_hd__xnor2_2 _29943_ (.A(_01383_),
    .B(_01391_),
    .Y(_01393_));
 sky130_fd_sc_hd__nand3_2 _29944_ (.A(_01380_),
    .B(_01382_),
    .C(_01393_),
    .Y(_01394_));
 sky130_fd_sc_hd__a21o_2 _29945_ (.A1(_01380_),
    .A2(_01382_),
    .B1(_01393_),
    .X(_01395_));
 sky130_fd_sc_hd__nand2_2 _29946_ (.A(_01394_),
    .B(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hd__nand2_2 _29947_ (.A(_01156_),
    .B(_01170_),
    .Y(_01397_));
 sky130_fd_sc_hd__xnor2_2 _29948_ (.A(_01396_),
    .B(_01397_),
    .Y(_01398_));
 sky130_fd_sc_hd__a21o_2 _29949_ (.A1(_01361_),
    .A2(_01362_),
    .B1(_01398_),
    .X(_01399_));
 sky130_fd_sc_hd__and3_2 _29950_ (.A(_01398_),
    .B(_01361_),
    .C(_01362_),
    .X(_01400_));
 sky130_fd_sc_hd__inv_2 _29951_ (.A(_01400_),
    .Y(_01401_));
 sky130_fd_sc_hd__o211ai_2 _29952_ (.A1(_01339_),
    .A2(_01200_),
    .B1(_01399_),
    .C1(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__a211o_2 _29953_ (.A1(_01399_),
    .A2(_01401_),
    .B1(_01339_),
    .C1(_01200_),
    .X(_01404_));
 sky130_fd_sc_hd__nand2_2 _29954_ (.A(_01402_),
    .B(_01404_),
    .Y(_01405_));
 sky130_fd_sc_hd__inv_2 _29955_ (.A(_01237_),
    .Y(_01406_));
 sky130_fd_sc_hd__and4_2 _29956_ (.A(iX[39]),
    .B(iX[40]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_01407_));
 sky130_fd_sc_hd__a22oi_2 _29957_ (.A1(iX[40]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[39]),
    .Y(_01408_));
 sky130_fd_sc_hd__nor2_2 _29958_ (.A(_01407_),
    .B(_01408_),
    .Y(_01409_));
 sky130_fd_sc_hd__nand2_2 _29959_ (.A(iX[38]),
    .B(iY[55]),
    .Y(_01410_));
 sky130_fd_sc_hd__xnor2_2 _29960_ (.A(_01409_),
    .B(_01410_),
    .Y(_01411_));
 sky130_fd_sc_hd__and4_2 _29961_ (.A(iX[42]),
    .B(iX[43]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_01412_));
 sky130_fd_sc_hd__a22oi_2 _29962_ (.A1(iX[43]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[42]),
    .Y(_01413_));
 sky130_fd_sc_hd__nor2_2 _29963_ (.A(_01412_),
    .B(_01413_),
    .Y(_01415_));
 sky130_fd_sc_hd__nand2_2 _29964_ (.A(iX[41]),
    .B(iY[52]),
    .Y(_01416_));
 sky130_fd_sc_hd__xnor2_2 _29965_ (.A(_01415_),
    .B(_01416_),
    .Y(_01417_));
 sky130_fd_sc_hd__o21ba_2 _29966_ (.A1(_01214_),
    .A2(_01216_),
    .B1_N(_01213_),
    .X(_01418_));
 sky130_fd_sc_hd__xnor2_2 _29967_ (.A(_01417_),
    .B(_01418_),
    .Y(_01419_));
 sky130_fd_sc_hd__and2_2 _29968_ (.A(_01411_),
    .B(_01419_),
    .X(_01420_));
 sky130_fd_sc_hd__nor2_2 _29969_ (.A(_01411_),
    .B(_01419_),
    .Y(_01421_));
 sky130_fd_sc_hd__or2_2 _29970_ (.A(_01420_),
    .B(_01421_),
    .X(_01422_));
 sky130_fd_sc_hd__or3_2 _29971_ (.A(_01225_),
    .B(_01230_),
    .C(_01231_),
    .X(_01423_));
 sky130_fd_sc_hd__o21ba_2 _29972_ (.A1(_01180_),
    .A2(_01182_),
    .B1_N(_01179_),
    .X(_01424_));
 sky130_fd_sc_hd__and4_2 _29973_ (.A(iX[45]),
    .B(iX[46]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_01426_));
 sky130_fd_sc_hd__a22oi_2 _29974_ (.A1(iX[46]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[45]),
    .Y(_01427_));
 sky130_fd_sc_hd__nand2_2 _29975_ (.A(iX[44]),
    .B(iY[49]),
    .Y(_01428_));
 sky130_fd_sc_hd__o21a_2 _29976_ (.A1(_01426_),
    .A2(_01427_),
    .B1(_01428_),
    .X(_01429_));
 sky130_fd_sc_hd__nor3_2 _29977_ (.A(_01426_),
    .B(_01427_),
    .C(_01428_),
    .Y(_01430_));
 sky130_fd_sc_hd__nor2_2 _29978_ (.A(_01429_),
    .B(_01430_),
    .Y(_01431_));
 sky130_fd_sc_hd__xnor2_2 _29979_ (.A(_01424_),
    .B(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__o21ai_2 _29980_ (.A1(_01226_),
    .A2(_01231_),
    .B1(_01432_),
    .Y(_01433_));
 sky130_fd_sc_hd__or3_2 _29981_ (.A(_01226_),
    .B(_01231_),
    .C(_01432_),
    .X(_01434_));
 sky130_fd_sc_hd__nand2_2 _29982_ (.A(_01433_),
    .B(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__a21oi_2 _29983_ (.A1(_01423_),
    .A2(_01234_),
    .B1(_01435_),
    .Y(_01437_));
 sky130_fd_sc_hd__and3_2 _29984_ (.A(_01423_),
    .B(_01234_),
    .C(_01435_),
    .X(_01438_));
 sky130_fd_sc_hd__or3_2 _29985_ (.A(_01422_),
    .B(_01437_),
    .C(_01438_),
    .X(_01439_));
 sky130_fd_sc_hd__o21ai_2 _29986_ (.A1(_01437_),
    .A2(_01438_),
    .B1(_01422_),
    .Y(_01440_));
 sky130_fd_sc_hd__nand2_2 _29987_ (.A(_01439_),
    .B(_01440_),
    .Y(_01441_));
 sky130_fd_sc_hd__a21oi_2 _29988_ (.A1(_01196_),
    .A2(_01198_),
    .B1(_01441_),
    .Y(_01442_));
 sky130_fd_sc_hd__and3_2 _29989_ (.A(_01196_),
    .B(_01198_),
    .C(_01441_),
    .X(_01443_));
 sky130_fd_sc_hd__a211oi_2 _29990_ (.A1(_01406_),
    .A2(_01240_),
    .B1(_01442_),
    .C1(_01443_),
    .Y(_01444_));
 sky130_fd_sc_hd__o211a_2 _29991_ (.A1(_01442_),
    .A2(_01443_),
    .B1(_01406_),
    .C1(_01240_),
    .X(_01445_));
 sky130_fd_sc_hd__or3_2 _29992_ (.A(_01405_),
    .B(_01444_),
    .C(_01445_),
    .X(_01446_));
 sky130_fd_sc_hd__inv_2 _29993_ (.A(_01446_),
    .Y(_01448_));
 sky130_fd_sc_hd__o21a_2 _29994_ (.A1(_01444_),
    .A2(_01445_),
    .B1(_01405_),
    .X(_01449_));
 sky130_fd_sc_hd__a211o_2 _29995_ (.A1(_01203_),
    .A2(_01247_),
    .B1(_01448_),
    .C1(_01449_),
    .X(_01450_));
 sky130_fd_sc_hd__inv_2 _29996_ (.A(_01450_),
    .Y(_01451_));
 sky130_fd_sc_hd__o211a_2 _29997_ (.A1(_01448_),
    .A2(_01449_),
    .B1(_01203_),
    .C1(_01247_),
    .X(_01452_));
 sky130_fd_sc_hd__nor2_2 _29998_ (.A(_01451_),
    .B(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__and4_2 _29999_ (.A(iX[33]),
    .B(iX[34]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_01454_));
 sky130_fd_sc_hd__a22oi_2 _30000_ (.A1(iX[34]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[33]),
    .Y(_01455_));
 sky130_fd_sc_hd__nor2_2 _30001_ (.A(_01454_),
    .B(_01455_),
    .Y(_01456_));
 sky130_fd_sc_hd__nand2_2 _30002_ (.A(iX[32]),
    .B(iY[61]),
    .Y(_01457_));
 sky130_fd_sc_hd__xnor2_2 _30003_ (.A(_01456_),
    .B(_01457_),
    .Y(_01459_));
 sky130_fd_sc_hd__nand2_2 _30004_ (.A(_01256_),
    .B(_01459_),
    .Y(_01460_));
 sky130_fd_sc_hd__or2_2 _30005_ (.A(_01256_),
    .B(_01459_),
    .X(_01461_));
 sky130_fd_sc_hd__nand2_2 _30006_ (.A(_01460_),
    .B(_01461_),
    .Y(_01462_));
 sky130_fd_sc_hd__or2b_2 _30007_ (.A(_01263_),
    .B_N(_01268_),
    .X(_01463_));
 sky130_fd_sc_hd__or2b_2 _30008_ (.A(_01262_),
    .B_N(_01269_),
    .X(_01464_));
 sky130_fd_sc_hd__and2b_2 _30009_ (.A_N(_01219_),
    .B(_01218_),
    .X(_01465_));
 sky130_fd_sc_hd__o21ba_2 _30010_ (.A1(_01265_),
    .A2(_01267_),
    .B1_N(_01264_),
    .X(_01466_));
 sky130_fd_sc_hd__o21ba_2 _30011_ (.A1(_01209_),
    .A2(_01211_),
    .B1_N(_01208_),
    .X(_01467_));
 sky130_fd_sc_hd__and4_2 _30012_ (.A(iX[36]),
    .B(iX[37]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_01468_));
 sky130_fd_sc_hd__a22oi_2 _30013_ (.A1(iX[37]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[36]),
    .Y(_01470_));
 sky130_fd_sc_hd__nor2_2 _30014_ (.A(_01468_),
    .B(_01470_),
    .Y(_01471_));
 sky130_fd_sc_hd__nand2_2 _30015_ (.A(iX[35]),
    .B(iY[58]),
    .Y(_01472_));
 sky130_fd_sc_hd__xnor2_2 _30016_ (.A(_01471_),
    .B(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__xnor2_2 _30017_ (.A(_01467_),
    .B(_01473_),
    .Y(_01474_));
 sky130_fd_sc_hd__xnor2_2 _30018_ (.A(_01466_),
    .B(_01474_),
    .Y(_01475_));
 sky130_fd_sc_hd__o21a_2 _30019_ (.A1(_01465_),
    .A2(_01221_),
    .B1(_01475_),
    .X(_01476_));
 sky130_fd_sc_hd__nor3_2 _30020_ (.A(_01465_),
    .B(_01221_),
    .C(_01475_),
    .Y(_01477_));
 sky130_fd_sc_hd__a211oi_2 _30021_ (.A1(_01463_),
    .A2(_01464_),
    .B1(_01476_),
    .C1(_01477_),
    .Y(_01478_));
 sky130_fd_sc_hd__o211a_2 _30022_ (.A1(_01476_),
    .A2(_01477_),
    .B1(_01463_),
    .C1(_01464_),
    .X(_01479_));
 sky130_fd_sc_hd__nor2_2 _30023_ (.A(_01478_),
    .B(_01479_),
    .Y(_01481_));
 sky130_fd_sc_hd__o21a_2 _30024_ (.A1(_01271_),
    .A2(_01274_),
    .B1(_01481_),
    .X(_01482_));
 sky130_fd_sc_hd__nor3_2 _30025_ (.A(_01271_),
    .B(_01274_),
    .C(_01481_),
    .Y(_01483_));
 sky130_fd_sc_hd__or3_2 _30026_ (.A(_01462_),
    .B(_01482_),
    .C(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__o21ai_2 _30027_ (.A1(_01482_),
    .A2(_01483_),
    .B1(_01462_),
    .Y(_01485_));
 sky130_fd_sc_hd__o211a_2 _30028_ (.A1(_01243_),
    .A2(_01245_),
    .B1(_01484_),
    .C1(_01485_),
    .X(_01486_));
 sky130_fd_sc_hd__a211oi_2 _30029_ (.A1(_01484_),
    .A2(_01485_),
    .B1(_01243_),
    .C1(_01245_),
    .Y(_01487_));
 sky130_fd_sc_hd__a211oi_2 _30030_ (.A1(_01277_),
    .A2(_01279_),
    .B1(_01486_),
    .C1(_01487_),
    .Y(_01488_));
 sky130_fd_sc_hd__o211a_2 _30031_ (.A1(_01486_),
    .A2(_01487_),
    .B1(_01277_),
    .C1(_01279_),
    .X(_01489_));
 sky130_fd_sc_hd__nor2_2 _30032_ (.A(_01488_),
    .B(_01489_),
    .Y(_01490_));
 sky130_fd_sc_hd__xnor2_2 _30033_ (.A(_01453_),
    .B(_01490_),
    .Y(_01492_));
 sky130_fd_sc_hd__a21o_2 _30034_ (.A1(_01254_),
    .A2(_01286_),
    .B1(_01252_),
    .X(_01493_));
 sky130_fd_sc_hd__xnor2_2 _30035_ (.A(_01492_),
    .B(_01493_),
    .Y(_01494_));
 sky130_fd_sc_hd__nor2_2 _30036_ (.A(_01281_),
    .B(_01284_),
    .Y(_01495_));
 sky130_fd_sc_hd__xnor2_2 _30037_ (.A(_01494_),
    .B(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__o21a_2 _30038_ (.A1(_01288_),
    .A2(_01290_),
    .B1(_01496_),
    .X(_01497_));
 sky130_fd_sc_hd__nor3_2 _30039_ (.A(_01288_),
    .B(_01290_),
    .C(_01496_),
    .Y(_01498_));
 sky130_fd_sc_hd__nor2_2 _30040_ (.A(_01497_),
    .B(_01498_),
    .Y(_01499_));
 sky130_fd_sc_hd__nand2_2 _30041_ (.A(_01338_),
    .B(_01499_),
    .Y(_01500_));
 sky130_fd_sc_hd__or2_2 _30042_ (.A(_01338_),
    .B(_01499_),
    .X(_01501_));
 sky130_fd_sc_hd__and2_2 _30043_ (.A(_01500_),
    .B(_01501_),
    .X(_01503_));
 sky130_fd_sc_hd__and2b_2 _30044_ (.A_N(_00871_),
    .B(_01295_),
    .X(_01504_));
 sky130_fd_sc_hd__nor2_2 _30045_ (.A(_01504_),
    .B(_01297_),
    .Y(_01505_));
 sky130_fd_sc_hd__xnor2_2 _30046_ (.A(_01503_),
    .B(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__inv_2 _30047_ (.A(_00973_),
    .Y(_01507_));
 sky130_fd_sc_hd__o211a_2 _30048_ (.A1(_00696_),
    .A2(_00698_),
    .B1(_01109_),
    .C1(_01110_),
    .X(_01508_));
 sky130_fd_sc_hd__a211o_2 _30049_ (.A1(_00551_),
    .A2(_00949_),
    .B1(_00967_),
    .C1(_00968_),
    .X(_01509_));
 sky130_fd_sc_hd__nor2_2 _30050_ (.A(_00940_),
    .B(_00941_),
    .Y(_01510_));
 sky130_fd_sc_hd__nand2_2 _30051_ (.A(_15616_),
    .B(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__xnor2_2 _30052_ (.A(_00562_),
    .B(_00563_),
    .Y(_01512_));
 sky130_fd_sc_hd__nor2_2 _30053_ (.A(_16625_),
    .B(_01512_),
    .Y(_01514_));
 sky130_fd_sc_hd__a21oi_2 _30054_ (.A1(_17392_),
    .A2(_01510_),
    .B1(_01514_),
    .Y(_01515_));
 sky130_fd_sc_hd__o21ba_2 _30055_ (.A1(_00945_),
    .A2(_01511_),
    .B1_N(_01515_),
    .X(_01516_));
 sky130_fd_sc_hd__and2_2 _30056_ (.A(iY[29]),
    .B(iY[61]),
    .X(_01517_));
 sky130_fd_sc_hd__nor2_2 _30057_ (.A(iY[29]),
    .B(iY[61]),
    .Y(_01518_));
 sky130_fd_sc_hd__or2_2 _30058_ (.A(_01517_),
    .B(_01518_),
    .X(_01519_));
 sky130_fd_sc_hd__nor2_2 _30059_ (.A(_00937_),
    .B(_00940_),
    .Y(_01520_));
 sky130_fd_sc_hd__xor2_2 _30060_ (.A(_01519_),
    .B(_01520_),
    .X(_01521_));
 sky130_fd_sc_hd__buf_1 _30061_ (.A(_01521_),
    .X(_01522_));
 sky130_fd_sc_hd__nand2_2 _30062_ (.A(_14592_),
    .B(_01522_),
    .Y(_01523_));
 sky130_fd_sc_hd__xor2_2 _30063_ (.A(_01516_),
    .B(_01523_),
    .X(_01525_));
 sky130_fd_sc_hd__or2_2 _30064_ (.A(_00947_),
    .B(_01525_),
    .X(_01526_));
 sky130_fd_sc_hd__nand2_2 _30065_ (.A(_00947_),
    .B(_01525_),
    .Y(_01527_));
 sky130_fd_sc_hd__and2_2 _30066_ (.A(_01526_),
    .B(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__nand3_2 _30067_ (.A(_00950_),
    .B(_00965_),
    .C(_00966_),
    .Y(_01529_));
 sky130_fd_sc_hd__nand2_2 _30068_ (.A(_00960_),
    .B(_00962_),
    .Y(_01530_));
 sky130_fd_sc_hd__nor2_2 _30069_ (.A(_00992_),
    .B(_00993_),
    .Y(_01531_));
 sky130_fd_sc_hd__a21o_2 _30070_ (.A1(_00984_),
    .A2(_00994_),
    .B1(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__nand2_2 _30071_ (.A(_00956_),
    .B(_00959_),
    .Y(_01533_));
 sky130_fd_sc_hd__o21bai_2 _30072_ (.A1(_00980_),
    .A2(_00981_),
    .B1_N(_00979_),
    .Y(_01534_));
 sky130_fd_sc_hd__or4b_2 _30073_ (.A(_14346_),
    .B(_14640_),
    .C(_18342_),
    .D_N(_18728_),
    .X(_01536_));
 sky130_fd_sc_hd__a22o_2 _30074_ (.A1(_15624_),
    .A2(_18732_),
    .B1(_18728_),
    .B2(_14628_),
    .X(_01537_));
 sky130_fd_sc_hd__a22o_2 _30075_ (.A1(_18749_),
    .A2(_00161_),
    .B1(_01536_),
    .B2(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__nand4_2 _30076_ (.A(_18749_),
    .B(_00162_),
    .C(_01536_),
    .D(_01537_),
    .Y(_01539_));
 sky130_fd_sc_hd__nand3_2 _30077_ (.A(_01534_),
    .B(_01538_),
    .C(_01539_),
    .Y(_01540_));
 sky130_fd_sc_hd__a21o_2 _30078_ (.A1(_01538_),
    .A2(_01539_),
    .B1(_01534_),
    .X(_01541_));
 sky130_fd_sc_hd__nand3_2 _30079_ (.A(_01533_),
    .B(_01540_),
    .C(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__a21o_2 _30080_ (.A1(_01540_),
    .A2(_01541_),
    .B1(_01533_),
    .X(_01543_));
 sky130_fd_sc_hd__nand3_2 _30081_ (.A(_01532_),
    .B(_01542_),
    .C(_01543_),
    .Y(_01544_));
 sky130_fd_sc_hd__a21o_2 _30082_ (.A1(_01542_),
    .A2(_01543_),
    .B1(_01532_),
    .X(_01545_));
 sky130_fd_sc_hd__and3_2 _30083_ (.A(_01530_),
    .B(_01544_),
    .C(_01545_),
    .X(_01547_));
 sky130_fd_sc_hd__a21oi_2 _30084_ (.A1(_01544_),
    .A2(_01545_),
    .B1(_01530_),
    .Y(_01548_));
 sky130_fd_sc_hd__a211o_2 _30085_ (.A1(_00965_),
    .A2(_01529_),
    .B1(_01547_),
    .C1(_01548_),
    .X(_01549_));
 sky130_fd_sc_hd__o211ai_2 _30086_ (.A1(_01547_),
    .A2(_01548_),
    .B1(_00965_),
    .C1(_01529_),
    .Y(_01550_));
 sky130_fd_sc_hd__and3_2 _30087_ (.A(_01528_),
    .B(_01549_),
    .C(_01550_),
    .X(_01551_));
 sky130_fd_sc_hd__a21oi_2 _30088_ (.A1(_01549_),
    .A2(_01550_),
    .B1(_01528_),
    .Y(_01552_));
 sky130_fd_sc_hd__a211oi_2 _30089_ (.A1(_01018_),
    .A2(_01021_),
    .B1(_01551_),
    .C1(_01552_),
    .Y(_01553_));
 sky130_fd_sc_hd__o211a_2 _30090_ (.A1(_01551_),
    .A2(_01552_),
    .B1(_01018_),
    .C1(_01021_),
    .X(_01554_));
 sky130_fd_sc_hd__a211oi_2 _30091_ (.A1(_01509_),
    .A2(_00971_),
    .B1(_01553_),
    .C1(_01554_),
    .Y(_01555_));
 sky130_fd_sc_hd__o211a_2 _30092_ (.A1(_01553_),
    .A2(_01554_),
    .B1(_01509_),
    .C1(_00971_),
    .X(_01556_));
 sky130_fd_sc_hd__nand2_2 _30093_ (.A(_00995_),
    .B(_01016_),
    .Y(_01558_));
 sky130_fd_sc_hd__and2b_2 _30094_ (.A_N(_01027_),
    .B(_01048_),
    .X(_01559_));
 sky130_fd_sc_hd__and2b_2 _30095_ (.A_N(_01025_),
    .B(_01049_),
    .X(_01560_));
 sky130_fd_sc_hd__and4_2 _30096_ (.A(_16277_),
    .B(_14652_),
    .C(_17630_),
    .D(_18101_),
    .X(_01561_));
 sky130_fd_sc_hd__a22o_2 _30097_ (.A1(_14652_),
    .A2(_17630_),
    .B1(_18101_),
    .B2(_16277_),
    .X(_01562_));
 sky130_fd_sc_hd__and2b_2 _30098_ (.A_N(_01561_),
    .B(_01562_),
    .X(_01563_));
 sky130_fd_sc_hd__buf_1 _30099_ (.A(_16268_),
    .X(_01564_));
 sky130_fd_sc_hd__nand2_2 _30100_ (.A(_01564_),
    .B(_18328_),
    .Y(_01565_));
 sky130_fd_sc_hd__xnor2_2 _30101_ (.A(_01563_),
    .B(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__or3b_2 _30102_ (.A(_15648_),
    .B(_16617_),
    .C_N(_00985_),
    .X(_01567_));
 sky130_fd_sc_hd__a2bb2o_2 _30103_ (.A1_N(_15648_),
    .A2_N(_16257_),
    .B1(_16614_),
    .B2(_00999_),
    .X(_01569_));
 sky130_fd_sc_hd__nand2_2 _30104_ (.A(_01567_),
    .B(_01569_),
    .Y(_01570_));
 sky130_fd_sc_hd__or2_2 _30105_ (.A(_16288_),
    .B(_18363_),
    .X(_01571_));
 sky130_fd_sc_hd__xnor2_2 _30106_ (.A(_01570_),
    .B(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__o21a_2 _30107_ (.A1(_00989_),
    .A2(_00991_),
    .B1(_00987_),
    .X(_01573_));
 sky130_fd_sc_hd__xor2_2 _30108_ (.A(_01572_),
    .B(_01573_),
    .X(_01574_));
 sky130_fd_sc_hd__xor2_2 _30109_ (.A(_01566_),
    .B(_01574_),
    .X(_01575_));
 sky130_fd_sc_hd__buf_1 _30110_ (.A(_15648_),
    .X(_01576_));
 sky130_fd_sc_hd__o31a_2 _30111_ (.A1(_01576_),
    .A2(_00996_),
    .A3(_01005_),
    .B1(_01003_),
    .X(_01577_));
 sky130_fd_sc_hd__or3_2 _30112_ (.A(_15169_),
    .B(_18181_),
    .C(_01029_),
    .X(_01578_));
 sky130_fd_sc_hd__o21a_2 _30113_ (.A1(_01031_),
    .A2(_01034_),
    .B1(_01578_),
    .X(_01580_));
 sky130_fd_sc_hd__nor2_2 _30114_ (.A(_14998_),
    .B(_15154_),
    .Y(_01581_));
 sky130_fd_sc_hd__xnor2_2 _30115_ (.A(_01002_),
    .B(_01581_),
    .Y(_01582_));
 sky130_fd_sc_hd__buf_1 _30116_ (.A(_14988_),
    .X(_01583_));
 sky130_fd_sc_hd__nor2_2 _30117_ (.A(_01583_),
    .B(_15835_),
    .Y(_01584_));
 sky130_fd_sc_hd__xnor2_2 _30118_ (.A(_01582_),
    .B(_01584_),
    .Y(_01585_));
 sky130_fd_sc_hd__xnor2_2 _30119_ (.A(_01580_),
    .B(_01585_),
    .Y(_01586_));
 sky130_fd_sc_hd__xnor2_2 _30120_ (.A(_01577_),
    .B(_01586_),
    .Y(_01587_));
 sky130_fd_sc_hd__and2b_2 _30121_ (.A_N(_01001_),
    .B(_01007_),
    .X(_01588_));
 sky130_fd_sc_hd__a21oi_2 _30122_ (.A1(_01000_),
    .A2(_01009_),
    .B1(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__xnor2_2 _30123_ (.A(_01587_),
    .B(_01589_),
    .Y(_01591_));
 sky130_fd_sc_hd__nand2_2 _30124_ (.A(_01575_),
    .B(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__or2_2 _30125_ (.A(_01575_),
    .B(_01591_),
    .X(_01593_));
 sky130_fd_sc_hd__o211a_2 _30126_ (.A1(_01559_),
    .A2(_01560_),
    .B1(_01592_),
    .C1(_01593_),
    .X(_01594_));
 sky130_fd_sc_hd__a211oi_2 _30127_ (.A1(_01592_),
    .A2(_01593_),
    .B1(_01559_),
    .C1(_01560_),
    .Y(_01595_));
 sky130_fd_sc_hd__a211oi_2 _30128_ (.A1(_01013_),
    .A2(_01558_),
    .B1(_01594_),
    .C1(_01595_),
    .Y(_01596_));
 sky130_fd_sc_hd__o211a_2 _30129_ (.A1(_01594_),
    .A2(_01595_),
    .B1(_01013_),
    .C1(_01558_),
    .X(_01597_));
 sky130_fd_sc_hd__inv_2 _30130_ (.A(_01102_),
    .Y(_01598_));
 sky130_fd_sc_hd__o21ai_2 _30131_ (.A1(_01035_),
    .A2(_01047_),
    .B1(_01045_),
    .Y(_01599_));
 sky130_fd_sc_hd__and2b_2 _30132_ (.A_N(_01060_),
    .B(_01054_),
    .X(_01600_));
 sky130_fd_sc_hd__and2b_2 _30133_ (.A_N(_01061_),
    .B(_01053_),
    .X(_01602_));
 sky130_fd_sc_hd__or2_2 _30134_ (.A(_01600_),
    .B(_01602_),
    .X(_01603_));
 sky130_fd_sc_hd__and3b_2 _30135_ (.A_N(_01029_),
    .B(_14608_),
    .C(_15900_),
    .X(_01604_));
 sky130_fd_sc_hd__buf_1 _30136_ (.A(_15168_),
    .X(_01605_));
 sky130_fd_sc_hd__o22a_2 _30137_ (.A1(_15169_),
    .A2(_16312_),
    .B1(_17696_),
    .B2(_01605_),
    .X(_01606_));
 sky130_fd_sc_hd__nor2_2 _30138_ (.A(_01604_),
    .B(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__a21oi_2 _30139_ (.A1(_01033_),
    .A2(_17460_),
    .B1(_01607_),
    .Y(_01608_));
 sky130_fd_sc_hd__and3_2 _30140_ (.A(_01033_),
    .B(_17460_),
    .C(_01607_),
    .X(_01609_));
 sky130_fd_sc_hd__or2_2 _30141_ (.A(_01608_),
    .B(_01609_),
    .X(_01610_));
 sky130_fd_sc_hd__nor2_2 _30142_ (.A(_13893_),
    .B(_01058_),
    .Y(_01611_));
 sky130_fd_sc_hd__o22a_2 _30143_ (.A1(_13893_),
    .A2(_17007_),
    .B1(_16999_),
    .B2(_14612_),
    .X(_01613_));
 sky130_fd_sc_hd__a21o_2 _30144_ (.A1(_01037_),
    .A2(_01611_),
    .B1(_01613_),
    .X(_01614_));
 sky130_fd_sc_hd__nand2_2 _30145_ (.A(_01039_),
    .B(_17006_),
    .Y(_01615_));
 sky130_fd_sc_hd__xnor2_2 _30146_ (.A(_01614_),
    .B(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__nand2_2 _30147_ (.A(_01036_),
    .B(_01037_),
    .Y(_01617_));
 sky130_fd_sc_hd__o21a_2 _30148_ (.A1(_01038_),
    .A2(_01042_),
    .B1(_01617_),
    .X(_01618_));
 sky130_fd_sc_hd__or2_2 _30149_ (.A(_01616_),
    .B(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__nand2_2 _30150_ (.A(_01616_),
    .B(_01618_),
    .Y(_01620_));
 sky130_fd_sc_hd__nand2_2 _30151_ (.A(_01619_),
    .B(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__xor2_2 _30152_ (.A(_01610_),
    .B(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__xnor2_2 _30153_ (.A(_01603_),
    .B(_01622_),
    .Y(_01624_));
 sky130_fd_sc_hd__xnor2_2 _30154_ (.A(_01599_),
    .B(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__inv_2 _30155_ (.A(_01098_),
    .Y(_01626_));
 sky130_fd_sc_hd__nor2_2 _30156_ (.A(_01058_),
    .B(_01057_),
    .Y(_01627_));
 sky130_fd_sc_hd__a22o_2 _30157_ (.A1(_01055_),
    .A2(_01056_),
    .B1(_01627_),
    .B2(_17463_),
    .X(_01628_));
 sky130_fd_sc_hd__or3b_2 _30158_ (.A(_14978_),
    .B(_00666_),
    .C_N(_00659_),
    .X(_01629_));
 sky130_fd_sc_hd__o31ai_2 _30159_ (.A1(_15646_),
    .A2(_01066_),
    .A3(_01064_),
    .B1(_01629_),
    .Y(_01630_));
 sky130_fd_sc_hd__nor2_2 _30160_ (.A(_14626_),
    .B(_18200_),
    .Y(_01631_));
 sky130_fd_sc_hd__or3b_2 _30161_ (.A(_12852_),
    .B(_18211_),
    .C_N(_01056_),
    .X(_01632_));
 sky130_fd_sc_hd__a22o_2 _30162_ (.A1(_14637_),
    .A2(_18463_),
    .B1(_00662_),
    .B2(_14636_),
    .X(_01633_));
 sky130_fd_sc_hd__nand3_2 _30163_ (.A(_01631_),
    .B(_01632_),
    .C(_01633_),
    .Y(_01635_));
 sky130_fd_sc_hd__a21o_2 _30164_ (.A1(_01632_),
    .A2(_01633_),
    .B1(_01631_),
    .X(_01636_));
 sky130_fd_sc_hd__nand3_2 _30165_ (.A(_01630_),
    .B(_01635_),
    .C(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__a21o_2 _30166_ (.A1(_01635_),
    .A2(_01636_),
    .B1(_01630_),
    .X(_01638_));
 sky130_fd_sc_hd__and3_2 _30167_ (.A(_01628_),
    .B(_01637_),
    .C(_01638_),
    .X(_01639_));
 sky130_fd_sc_hd__a21oi_2 _30168_ (.A1(_01637_),
    .A2(_01638_),
    .B1(_01628_),
    .Y(_01640_));
 sky130_fd_sc_hd__nor2_2 _30169_ (.A(_01639_),
    .B(_01640_),
    .Y(_01641_));
 sky130_fd_sc_hd__nand2_2 _30170_ (.A(_14980_),
    .B(_00268_),
    .Y(_01642_));
 sky130_fd_sc_hd__nor2_2 _30171_ (.A(_00278_),
    .B(_00280_),
    .Y(_01643_));
 sky130_fd_sc_hd__nand2_2 _30172_ (.A(_14649_),
    .B(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__xor2_2 _30173_ (.A(_01642_),
    .B(_01644_),
    .X(_01646_));
 sky130_fd_sc_hd__buf_1 _30174_ (.A(_18460_),
    .X(_01647_));
 sky130_fd_sc_hd__nand2_2 _30175_ (.A(_18192_),
    .B(_01647_),
    .Y(_01648_));
 sky130_fd_sc_hd__xnor2_2 _30176_ (.A(_01646_),
    .B(_01648_),
    .Y(_01649_));
 sky130_fd_sc_hd__nor2_2 _30177_ (.A(_00674_),
    .B(_00675_),
    .Y(_01650_));
 sky130_fd_sc_hd__a21o_2 _30178_ (.A1(_01075_),
    .A2(_01077_),
    .B1(_01080_),
    .X(_01651_));
 sky130_fd_sc_hd__or2_2 _30179_ (.A(iX[29]),
    .B(iX[61]),
    .X(_01652_));
 sky130_fd_sc_hd__nand2_2 _30180_ (.A(iX[29]),
    .B(iX[61]),
    .Y(_01653_));
 sky130_fd_sc_hd__nand2_2 _30181_ (.A(_01652_),
    .B(_01653_),
    .Y(_01654_));
 sky130_fd_sc_hd__and3_2 _30182_ (.A(_01078_),
    .B(_01651_),
    .C(_01654_),
    .X(_01655_));
 sky130_fd_sc_hd__a21oi_2 _30183_ (.A1(_01078_),
    .A2(_01651_),
    .B1(_01654_),
    .Y(_01657_));
 sky130_fd_sc_hd__or4_2 _30184_ (.A(_11566_),
    .B(_01083_),
    .C(_01655_),
    .D(_01657_),
    .X(_01658_));
 sky130_fd_sc_hd__o31ai_2 _30185_ (.A1(_11567_),
    .A2(_01655_),
    .A3(_01657_),
    .B1(_01083_),
    .Y(_01659_));
 sky130_fd_sc_hd__nand4_2 _30186_ (.A(_15677_),
    .B(_01650_),
    .C(_01658_),
    .D(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__a22o_2 _30187_ (.A1(_15677_),
    .A2(_01650_),
    .B1(_01658_),
    .B2(_01659_),
    .X(_01661_));
 sky130_fd_sc_hd__a21bo_2 _30188_ (.A1(_01071_),
    .A2(_01088_),
    .B1_N(_01084_),
    .X(_01662_));
 sky130_fd_sc_hd__nand3_2 _30189_ (.A(_01660_),
    .B(_01661_),
    .C(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__a21o_2 _30190_ (.A1(_01660_),
    .A2(_01661_),
    .B1(_01662_),
    .X(_01664_));
 sky130_fd_sc_hd__nand3_2 _30191_ (.A(_01649_),
    .B(_01663_),
    .C(_01664_),
    .Y(_01665_));
 sky130_fd_sc_hd__a21o_2 _30192_ (.A1(_01663_),
    .A2(_01664_),
    .B1(_01649_),
    .X(_01666_));
 sky130_fd_sc_hd__a21bo_2 _30193_ (.A1(_01068_),
    .A2(_01093_),
    .B1_N(_01092_),
    .X(_01668_));
 sky130_fd_sc_hd__nand3_2 _30194_ (.A(_01665_),
    .B(_01666_),
    .C(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__a21o_2 _30195_ (.A1(_01665_),
    .A2(_01666_),
    .B1(_01668_),
    .X(_01670_));
 sky130_fd_sc_hd__nand3_2 _30196_ (.A(_01641_),
    .B(_01669_),
    .C(_01670_),
    .Y(_01671_));
 sky130_fd_sc_hd__a21o_2 _30197_ (.A1(_01669_),
    .A2(_01670_),
    .B1(_01641_),
    .X(_01672_));
 sky130_fd_sc_hd__o211ai_2 _30198_ (.A1(_01626_),
    .A2(_01100_),
    .B1(_01671_),
    .C1(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hd__a211o_2 _30199_ (.A1(_01671_),
    .A2(_01672_),
    .B1(_01626_),
    .C1(_01100_),
    .X(_01674_));
 sky130_fd_sc_hd__nand3_2 _30200_ (.A(_01625_),
    .B(_01673_),
    .C(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__a21o_2 _30201_ (.A1(_01673_),
    .A2(_01674_),
    .B1(_01625_),
    .X(_01676_));
 sky130_fd_sc_hd__o211a_2 _30202_ (.A1(_01598_),
    .A2(_01104_),
    .B1(_01675_),
    .C1(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__a211oi_2 _30203_ (.A1(_01675_),
    .A2(_01676_),
    .B1(_01598_),
    .C1(_01104_),
    .Y(_01679_));
 sky130_fd_sc_hd__nor4_2 _30204_ (.A(_01596_),
    .B(_01597_),
    .C(_01677_),
    .D(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__o22a_2 _30205_ (.A1(_01596_),
    .A2(_01597_),
    .B1(_01677_),
    .B2(_01679_),
    .X(_01681_));
 sky130_fd_sc_hd__a211o_2 _30206_ (.A1(_01106_),
    .A2(_01109_),
    .B1(_01680_),
    .C1(_01681_),
    .X(_01682_));
 sky130_fd_sc_hd__o211ai_2 _30207_ (.A1(_01680_),
    .A2(_01681_),
    .B1(_01106_),
    .C1(_01109_),
    .Y(_01683_));
 sky130_fd_sc_hd__nand4bb_2 _30208_ (.A_N(_01555_),
    .B_N(_01556_),
    .C(_01682_),
    .D(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__a2bb2o_2 _30209_ (.A1_N(_01555_),
    .A2_N(_01556_),
    .B1(_01682_),
    .B2(_01683_),
    .X(_01685_));
 sky130_fd_sc_hd__o211a_2 _30210_ (.A1(_01508_),
    .A2(_01113_),
    .B1(_01684_),
    .C1(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__a211oi_2 _30211_ (.A1(_01684_),
    .A2(_01685_),
    .B1(_01508_),
    .C1(_01113_),
    .Y(_01687_));
 sky130_fd_sc_hd__a211oi_2 _30212_ (.A1(_01507_),
    .A2(_00976_),
    .B1(_01686_),
    .C1(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__o211a_2 _30213_ (.A1(_01686_),
    .A2(_01687_),
    .B1(_01507_),
    .C1(_00976_),
    .X(_01690_));
 sky130_fd_sc_hd__a211oi_2 _30214_ (.A1(_01115_),
    .A2(_01117_),
    .B1(_01688_),
    .C1(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__o211a_2 _30215_ (.A1(_01688_),
    .A2(_01690_),
    .B1(_01115_),
    .C1(_01117_),
    .X(_01692_));
 sky130_fd_sc_hd__o21a_2 _30216_ (.A1(_01691_),
    .A2(_01692_),
    .B1(_01120_),
    .X(_01693_));
 sky130_fd_sc_hd__or3_2 _30217_ (.A(_01120_),
    .B(_01691_),
    .C(_01692_),
    .X(_01694_));
 sky130_fd_sc_hd__or2b_2 _30218_ (.A(_01693_),
    .B_N(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__nor2_2 _30219_ (.A(_00709_),
    .B(_01122_),
    .Y(_01696_));
 sky130_fd_sc_hd__o21ba_2 _30220_ (.A1(_01123_),
    .A2(_01132_),
    .B1_N(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__xor2_2 _30221_ (.A(_01695_),
    .B(_01697_),
    .X(_01698_));
 sky130_fd_sc_hd__xnor2_2 _30222_ (.A(_01506_),
    .B(_01698_),
    .Y(_01699_));
 sky130_fd_sc_hd__xnor2_2 _30223_ (.A(_10830_),
    .B(_01699_),
    .Y(_01701_));
 sky130_fd_sc_hd__and3_2 _30224_ (.A(_01336_),
    .B(_01301_),
    .C(_01701_),
    .X(_01702_));
 sky130_fd_sc_hd__a21oi_2 _30225_ (.A1(_01336_),
    .A2(_01301_),
    .B1(_01701_),
    .Y(_01703_));
 sky130_fd_sc_hd__or2_2 _30226_ (.A(_01702_),
    .B(_01703_),
    .X(_01704_));
 sky130_fd_sc_hd__nor2_2 _30227_ (.A(_01303_),
    .B(_01304_),
    .Y(_01705_));
 sky130_fd_sc_hd__a311o_2 _30228_ (.A1(_00477_),
    .A2(_00479_),
    .A3(_00925_),
    .B1(_01306_),
    .C1(_00926_),
    .X(_01706_));
 sky130_fd_sc_hd__or2b_2 _30229_ (.A(_01705_),
    .B_N(_01706_),
    .X(_01707_));
 sky130_fd_sc_hd__xnor2_2 _30230_ (.A(_01704_),
    .B(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__nand2_2 _30231_ (.A(_01335_),
    .B(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__inv_2 _30232_ (.A(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hd__nor2_2 _30233_ (.A(_01335_),
    .B(_01708_),
    .Y(_01712_));
 sky130_fd_sc_hd__nor2_2 _30234_ (.A(_01710_),
    .B(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__inv_2 _30235_ (.A(_01310_),
    .Y(_01714_));
 sky130_fd_sc_hd__o221ai_2 _30236_ (.A1(_00097_),
    .A2(_01313_),
    .B1(_01314_),
    .B2(_01312_),
    .C1(_01714_),
    .Y(_01715_));
 sky130_fd_sc_hd__nand2_2 _30237_ (.A(_01308_),
    .B(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__xor2_2 _30238_ (.A(_01713_),
    .B(_01716_),
    .X(oO[61]));
 sky130_fd_sc_hd__or2b_2 _30239_ (.A(_00911_),
    .B_N(_01323_),
    .X(_01717_));
 sky130_fd_sc_hd__or2b_2 _30240_ (.A(_01325_),
    .B_N(_01324_),
    .X(_01718_));
 sky130_fd_sc_hd__nand2_2 _30241_ (.A(iX[31]),
    .B(iY[31]),
    .Y(_01719_));
 sky130_fd_sc_hd__o21ba_2 _30242_ (.A1(_01320_),
    .A2(_01322_),
    .B1_N(_01319_),
    .X(_01720_));
 sky130_fd_sc_hd__xnor2_2 _30243_ (.A(_01719_),
    .B(_01720_),
    .Y(_01722_));
 sky130_fd_sc_hd__a21o_2 _30244_ (.A1(_01717_),
    .A2(_01718_),
    .B1(_01722_),
    .X(_01723_));
 sky130_fd_sc_hd__nand3_2 _30245_ (.A(_01717_),
    .B(_01718_),
    .C(_01722_),
    .Y(_01724_));
 sky130_fd_sc_hd__nand2_2 _30246_ (.A(_01723_),
    .B(_01724_),
    .Y(_01725_));
 sky130_fd_sc_hd__o21ai_2 _30247_ (.A1(_01331_),
    .A2(_01333_),
    .B1(_01328_),
    .Y(_01726_));
 sky130_fd_sc_hd__or2b_2 _30248_ (.A(_01725_),
    .B_N(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__or2b_2 _30249_ (.A(_01726_),
    .B_N(_01725_),
    .X(_01728_));
 sky130_fd_sc_hd__nand2_2 _30250_ (.A(_01727_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__nor2_2 _30251_ (.A(_01705_),
    .B(_01703_),
    .Y(_01730_));
 sky130_fd_sc_hd__inv_2 _30252_ (.A(_01549_),
    .Y(_01731_));
 sky130_fd_sc_hd__buf_2 _30253_ (.A(_01510_),
    .X(_01733_));
 sky130_fd_sc_hd__o22a_2 _30254_ (.A1(_18120_),
    .A2(_01512_),
    .B1(_00943_),
    .B2(_16625_),
    .X(_01734_));
 sky130_fd_sc_hd__a31o_2 _30255_ (.A1(_18749_),
    .A2(_01733_),
    .A3(_01514_),
    .B1(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__nand2_2 _30256_ (.A(_17392_),
    .B(_01521_),
    .Y(_01736_));
 sky130_fd_sc_hd__xnor2_2 _30257_ (.A(_01735_),
    .B(_01736_),
    .Y(_01737_));
 sky130_fd_sc_hd__o22a_2 _30258_ (.A1(_00945_),
    .A2(_01511_),
    .B1(_01515_),
    .B2(_01523_),
    .X(_01738_));
 sky130_fd_sc_hd__xnor2_2 _30259_ (.A(_01737_),
    .B(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__nand2_2 _30260_ (.A(iY[30]),
    .B(iY[62]),
    .Y(_01740_));
 sky130_fd_sc_hd__or2_2 _30261_ (.A(iY[30]),
    .B(iY[62]),
    .X(_01741_));
 sky130_fd_sc_hd__nand2_2 _30262_ (.A(_01740_),
    .B(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__or2_2 _30263_ (.A(_00937_),
    .B(_01517_),
    .X(_01744_));
 sky130_fd_sc_hd__o21ba_2 _30264_ (.A1(_00940_),
    .A2(_01744_),
    .B1_N(_01518_),
    .X(_01745_));
 sky130_fd_sc_hd__xor2_2 _30265_ (.A(_01742_),
    .B(_01745_),
    .X(_01746_));
 sky130_fd_sc_hd__nor2_2 _30266_ (.A(_11579_),
    .B(_01746_),
    .Y(_01747_));
 sky130_fd_sc_hd__xnor2_2 _30267_ (.A(_01739_),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__xnor2_2 _30268_ (.A(_01526_),
    .B(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__nand3_2 _30269_ (.A(_01530_),
    .B(_01544_),
    .C(_01545_),
    .Y(_01750_));
 sky130_fd_sc_hd__nand2_2 _30270_ (.A(_01540_),
    .B(_01542_),
    .Y(_01751_));
 sky130_fd_sc_hd__nor2_2 _30271_ (.A(_01572_),
    .B(_01573_),
    .Y(_01752_));
 sky130_fd_sc_hd__a21o_2 _30272_ (.A1(_01566_),
    .A2(_01574_),
    .B1(_01752_),
    .X(_01753_));
 sky130_fd_sc_hd__nand2_2 _30273_ (.A(_01536_),
    .B(_01539_),
    .Y(_01755_));
 sky130_fd_sc_hd__a31o_2 _30274_ (.A1(_01564_),
    .A2(_18328_),
    .A3(_01562_),
    .B1(_01561_),
    .X(_01756_));
 sky130_fd_sc_hd__buf_6 _30275_ (.A(_00162_),
    .X(_01757_));
 sky130_fd_sc_hd__or4b_2 _30276_ (.A(_18368_),
    .B(_00195_),
    .C(_18343_),
    .D_N(_18728_),
    .X(_01758_));
 sky130_fd_sc_hd__a22o_2 _30277_ (.A1(_16268_),
    .A2(_18734_),
    .B1(_18729_),
    .B2(_18754_),
    .X(_01759_));
 sky130_fd_sc_hd__a22o_2 _30278_ (.A1(_14629_),
    .A2(_01757_),
    .B1(_01758_),
    .B2(_01759_),
    .X(_01760_));
 sky130_fd_sc_hd__nand4_2 _30279_ (.A(_14629_),
    .B(_01757_),
    .C(_01758_),
    .D(_01759_),
    .Y(_01761_));
 sky130_fd_sc_hd__nand3_2 _30280_ (.A(_01756_),
    .B(_01760_),
    .C(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__a21o_2 _30281_ (.A1(_01760_),
    .A2(_01761_),
    .B1(_01756_),
    .X(_01763_));
 sky130_fd_sc_hd__nand3_2 _30282_ (.A(_01755_),
    .B(_01762_),
    .C(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__a21o_2 _30283_ (.A1(_01762_),
    .A2(_01763_),
    .B1(_01755_),
    .X(_01766_));
 sky130_fd_sc_hd__nand3_2 _30284_ (.A(_01753_),
    .B(_01764_),
    .C(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__a21o_2 _30285_ (.A1(_01764_),
    .A2(_01766_),
    .B1(_01753_),
    .X(_01768_));
 sky130_fd_sc_hd__and3_4 _30286_ (.A(_01751_),
    .B(_01767_),
    .C(_01768_),
    .X(_01769_));
 sky130_fd_sc_hd__a21oi_2 _30287_ (.A1(_01767_),
    .A2(_01768_),
    .B1(_01751_),
    .Y(_01770_));
 sky130_fd_sc_hd__a211o_2 _30288_ (.A1(_01544_),
    .A2(_01750_),
    .B1(_01769_),
    .C1(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__o211ai_2 _30289_ (.A1(_01769_),
    .A2(_01770_),
    .B1(_01544_),
    .C1(_01750_),
    .Y(_01772_));
 sky130_fd_sc_hd__nand3_2 _30290_ (.A(_01749_),
    .B(_01771_),
    .C(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__a21o_2 _30291_ (.A1(_01771_),
    .A2(_01772_),
    .B1(_01749_),
    .X(_01774_));
 sky130_fd_sc_hd__o211ai_2 _30292_ (.A1(_01594_),
    .A2(_01596_),
    .B1(_01773_),
    .C1(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__a211o_2 _30293_ (.A1(_01773_),
    .A2(_01774_),
    .B1(_01594_),
    .C1(_01596_),
    .X(_01777_));
 sky130_fd_sc_hd__o211ai_2 _30294_ (.A1(_01731_),
    .A2(_01551_),
    .B1(_01775_),
    .C1(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__a211o_2 _30295_ (.A1(_01775_),
    .A2(_01777_),
    .B1(_01731_),
    .C1(_01551_),
    .X(_01779_));
 sky130_fd_sc_hd__or2b_2 _30296_ (.A(_01589_),
    .B_N(_01587_),
    .X(_01780_));
 sky130_fd_sc_hd__nand2_2 _30297_ (.A(_01780_),
    .B(_01592_),
    .Y(_01781_));
 sky130_fd_sc_hd__or2b_2 _30298_ (.A(_01624_),
    .B_N(_01599_),
    .X(_01782_));
 sky130_fd_sc_hd__a21bo_2 _30299_ (.A1(_01603_),
    .A2(_01622_),
    .B1_N(_01782_),
    .X(_01783_));
 sky130_fd_sc_hd__buf_1 _30300_ (.A(_14652_),
    .X(_01784_));
 sky130_fd_sc_hd__buf_1 _30301_ (.A(_14648_),
    .X(_01785_));
 sky130_fd_sc_hd__and4_2 _30302_ (.A(_01784_),
    .B(_01785_),
    .C(_17630_),
    .D(_18101_),
    .X(_01786_));
 sky130_fd_sc_hd__o22a_2 _30303_ (.A1(_16288_),
    .A2(_17408_),
    .B1(_17628_),
    .B2(_00990_),
    .X(_01788_));
 sky130_fd_sc_hd__or3_4 _30304_ (.A(_00589_),
    .B(_18111_),
    .C(_18113_),
    .X(_01789_));
 sky130_fd_sc_hd__o21a_2 _30305_ (.A1(_01786_),
    .A2(_01788_),
    .B1(_01789_),
    .X(_01790_));
 sky130_fd_sc_hd__or3_2 _30306_ (.A(_01786_),
    .B(_01788_),
    .C(_01789_),
    .X(_01791_));
 sky130_fd_sc_hd__nor2b_2 _30307_ (.A(_01790_),
    .B_N(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hd__nor2_2 _30308_ (.A(_14988_),
    .B(_16257_),
    .Y(_01793_));
 sky130_fd_sc_hd__or3b_2 _30309_ (.A(_15648_),
    .B(_16617_),
    .C_N(_01793_),
    .X(_01794_));
 sky130_fd_sc_hd__a21o_2 _30310_ (.A1(_18157_),
    .A2(_16614_),
    .B1(_01793_),
    .X(_01795_));
 sky130_fd_sc_hd__nand2_2 _30311_ (.A(_01794_),
    .B(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__buf_1 _30312_ (.A(_15211_),
    .X(_01797_));
 sky130_fd_sc_hd__or2_2 _30313_ (.A(_01797_),
    .B(_18363_),
    .X(_01799_));
 sky130_fd_sc_hd__xnor2_2 _30314_ (.A(_01796_),
    .B(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__o21a_2 _30315_ (.A1(_01570_),
    .A2(_01571_),
    .B1(_01567_),
    .X(_01801_));
 sky130_fd_sc_hd__xor2_2 _30316_ (.A(_01800_),
    .B(_01801_),
    .X(_01802_));
 sky130_fd_sc_hd__xor2_2 _30317_ (.A(_01792_),
    .B(_01802_),
    .X(_01803_));
 sky130_fd_sc_hd__buf_1 _30318_ (.A(_00996_),
    .X(_01804_));
 sky130_fd_sc_hd__nor2_2 _30319_ (.A(_01804_),
    .B(_01582_),
    .Y(_01805_));
 sky130_fd_sc_hd__a22o_2 _30320_ (.A1(_01002_),
    .A2(_01581_),
    .B1(_01805_),
    .B2(_15888_),
    .X(_01806_));
 sky130_fd_sc_hd__or2_2 _30321_ (.A(_14998_),
    .B(_15598_),
    .X(_01807_));
 sky130_fd_sc_hd__or3_2 _30322_ (.A(_15154_),
    .B(_15219_),
    .C(_15220_),
    .X(_01808_));
 sky130_fd_sc_hd__xnor2_2 _30323_ (.A(_01807_),
    .B(_01808_),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_2 _30324_ (.A(_15005_),
    .B(_00996_),
    .Y(_01811_));
 sky130_fd_sc_hd__xnor2_2 _30325_ (.A(_01810_),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__o21a_2 _30326_ (.A1(_01604_),
    .A2(_01609_),
    .B1(_01812_),
    .X(_01813_));
 sky130_fd_sc_hd__nor3_2 _30327_ (.A(_01604_),
    .B(_01609_),
    .C(_01812_),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_2 _30328_ (.A(_01813_),
    .B(_01814_),
    .Y(_01815_));
 sky130_fd_sc_hd__xor2_2 _30329_ (.A(_01806_),
    .B(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__and2b_2 _30330_ (.A_N(_01580_),
    .B(_01585_),
    .X(_01817_));
 sky130_fd_sc_hd__and2b_2 _30331_ (.A_N(_01577_),
    .B(_01586_),
    .X(_01818_));
 sky130_fd_sc_hd__nor2_2 _30332_ (.A(_01817_),
    .B(_01818_),
    .Y(_01819_));
 sky130_fd_sc_hd__xnor2_2 _30333_ (.A(_01816_),
    .B(_01819_),
    .Y(_01821_));
 sky130_fd_sc_hd__xnor2_2 _30334_ (.A(_01803_),
    .B(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__xor2_2 _30335_ (.A(_01783_),
    .B(_01822_),
    .X(_01823_));
 sky130_fd_sc_hd__xor2_2 _30336_ (.A(_01781_),
    .B(_01823_),
    .X(_01824_));
 sky130_fd_sc_hd__o21ai_2 _30337_ (.A1(_01610_),
    .A2(_01621_),
    .B1(_01619_),
    .Y(_01825_));
 sky130_fd_sc_hd__a31o_2 _30338_ (.A1(_01630_),
    .A2(_01635_),
    .A3(_01636_),
    .B1(_01639_),
    .X(_01826_));
 sky130_fd_sc_hd__and4_2 _30339_ (.A(_14411_),
    .B(_14606_),
    .C(_01040_),
    .D(_17006_),
    .X(_01827_));
 sky130_fd_sc_hd__buf_1 _30340_ (.A(_17696_),
    .X(_01828_));
 sky130_fd_sc_hd__o22a_2 _30341_ (.A1(_15169_),
    .A2(_01828_),
    .B1(_00255_),
    .B2(_01605_),
    .X(_01829_));
 sky130_fd_sc_hd__nor2_2 _30342_ (.A(_01827_),
    .B(_01829_),
    .Y(_01830_));
 sky130_fd_sc_hd__buf_1 _30343_ (.A(_16312_),
    .X(_01832_));
 sky130_fd_sc_hd__nor2_2 _30344_ (.A(_14949_),
    .B(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__xnor2_2 _30345_ (.A(_01830_),
    .B(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__nor2_2 _30346_ (.A(_18791_),
    .B(_17482_),
    .Y(_01835_));
 sky130_fd_sc_hd__xnor2_2 _30347_ (.A(_01611_),
    .B(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__buf_1 _30348_ (.A(_17488_),
    .X(_01837_));
 sky130_fd_sc_hd__nand2_2 _30349_ (.A(_01039_),
    .B(_01837_),
    .Y(_01838_));
 sky130_fd_sc_hd__xnor2_2 _30350_ (.A(_01836_),
    .B(_01838_),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_2 _30351_ (.A(_01037_),
    .B(_01611_),
    .Y(_01840_));
 sky130_fd_sc_hd__o21a_2 _30352_ (.A1(_01614_),
    .A2(_01615_),
    .B1(_01840_),
    .X(_01841_));
 sky130_fd_sc_hd__or2_2 _30353_ (.A(_01839_),
    .B(_01841_),
    .X(_01843_));
 sky130_fd_sc_hd__nand2_2 _30354_ (.A(_01839_),
    .B(_01841_),
    .Y(_01844_));
 sky130_fd_sc_hd__nand2_2 _30355_ (.A(_01843_),
    .B(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__xor2_2 _30356_ (.A(_01834_),
    .B(_01845_),
    .X(_01846_));
 sky130_fd_sc_hd__xnor2_2 _30357_ (.A(_01826_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__xnor2_2 _30358_ (.A(_01825_),
    .B(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__nor2_2 _30359_ (.A(_01642_),
    .B(_01644_),
    .Y(_01849_));
 sky130_fd_sc_hd__a31o_2 _30360_ (.A1(_18192_),
    .A2(_01647_),
    .A3(_01646_),
    .B1(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__nand2_2 _30361_ (.A(_17463_),
    .B(_18463_),
    .Y(_01851_));
 sky130_fd_sc_hd__nor2_2 _30362_ (.A(_12848_),
    .B(_18456_),
    .Y(_01852_));
 sky130_fd_sc_hd__or3b_2 _30363_ (.A(_12852_),
    .B(_18211_),
    .C_N(_01852_),
    .X(_01854_));
 sky130_fd_sc_hd__a21o_2 _30364_ (.A1(_14637_),
    .A2(_00662_),
    .B1(_01852_),
    .X(_01855_));
 sky130_fd_sc_hd__and2_2 _30365_ (.A(_01854_),
    .B(_01855_),
    .X(_01856_));
 sky130_fd_sc_hd__xnor2_2 _30366_ (.A(_01851_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__xnor2_2 _30367_ (.A(_01850_),
    .B(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__a21oi_2 _30368_ (.A1(_01632_),
    .A2(_01635_),
    .B1(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__and3_2 _30369_ (.A(_01632_),
    .B(_01635_),
    .C(_01858_),
    .X(_01860_));
 sky130_fd_sc_hd__or2_2 _30370_ (.A(_01859_),
    .B(_01860_),
    .X(_01861_));
 sky130_fd_sc_hd__buf_1 _30371_ (.A(_00268_),
    .X(_01862_));
 sky130_fd_sc_hd__nand2_2 _30372_ (.A(_18192_),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__or2_2 _30373_ (.A(_00674_),
    .B(_00675_),
    .X(_01865_));
 sky130_fd_sc_hd__buf_1 _30374_ (.A(_01865_),
    .X(_01866_));
 sky130_fd_sc_hd__nor3_2 _30375_ (.A(_14978_),
    .B(_01866_),
    .C(_01644_),
    .Y(_01867_));
 sky130_fd_sc_hd__a22o_2 _30376_ (.A1(_00661_),
    .A2(_01643_),
    .B1(_01650_),
    .B2(_14649_),
    .X(_01868_));
 sky130_fd_sc_hd__and2b_2 _30377_ (.A_N(_01867_),
    .B(_01868_),
    .X(_01869_));
 sky130_fd_sc_hd__xnor2_2 _30378_ (.A(_01863_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__nor2_2 _30379_ (.A(_11794_),
    .B(_01087_),
    .Y(_01871_));
 sky130_fd_sc_hd__or3_2 _30380_ (.A(_11576_),
    .B(_01655_),
    .C(_01657_),
    .X(_01872_));
 sky130_fd_sc_hd__and3_2 _30381_ (.A(iX[28]),
    .B(iX[60]),
    .C(_01652_),
    .X(_01873_));
 sky130_fd_sc_hd__a21oi_2 _30382_ (.A1(iX[29]),
    .A2(iX[61]),
    .B1(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__a211o_2 _30383_ (.A1(_01075_),
    .A2(_01077_),
    .B1(_01654_),
    .C1(_01080_),
    .X(_01876_));
 sky130_fd_sc_hd__nand2_2 _30384_ (.A(iX[30]),
    .B(iX[62]),
    .Y(_01877_));
 sky130_fd_sc_hd__or2_2 _30385_ (.A(iX[30]),
    .B(iX[62]),
    .X(_01878_));
 sky130_fd_sc_hd__nand2_2 _30386_ (.A(_01877_),
    .B(_01878_),
    .Y(_01879_));
 sky130_fd_sc_hd__a21o_2 _30387_ (.A1(_01874_),
    .A2(_01876_),
    .B1(_01879_),
    .X(_01880_));
 sky130_fd_sc_hd__nand3_2 _30388_ (.A(_01879_),
    .B(_01874_),
    .C(_01876_),
    .Y(_01881_));
 sky130_fd_sc_hd__and3_2 _30389_ (.A(_11381_),
    .B(_01880_),
    .C(_01881_),
    .X(_01882_));
 sky130_fd_sc_hd__xnor2_2 _30390_ (.A(_01872_),
    .B(_01882_),
    .Y(_01883_));
 sky130_fd_sc_hd__xnor2_2 _30391_ (.A(_01871_),
    .B(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__and2_2 _30392_ (.A(_01658_),
    .B(_01660_),
    .X(_01885_));
 sky130_fd_sc_hd__xor2_2 _30393_ (.A(_01884_),
    .B(_01885_),
    .X(_01887_));
 sky130_fd_sc_hd__xnor2_2 _30394_ (.A(_01870_),
    .B(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__and2_2 _30395_ (.A(_01663_),
    .B(_01665_),
    .X(_01889_));
 sky130_fd_sc_hd__xnor2_2 _30396_ (.A(_01888_),
    .B(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hd__xnor2_2 _30397_ (.A(_01861_),
    .B(_01890_),
    .Y(_01891_));
 sky130_fd_sc_hd__and2_2 _30398_ (.A(_01669_),
    .B(_01671_),
    .X(_01892_));
 sky130_fd_sc_hd__xor2_2 _30399_ (.A(_01891_),
    .B(_01892_),
    .X(_01893_));
 sky130_fd_sc_hd__xnor2_2 _30400_ (.A(_01848_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__and2_2 _30401_ (.A(_01673_),
    .B(_01675_),
    .X(_01895_));
 sky130_fd_sc_hd__xnor2_2 _30402_ (.A(_01894_),
    .B(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__xor2_2 _30403_ (.A(_01824_),
    .B(_01896_),
    .X(_01898_));
 sky130_fd_sc_hd__nor2_2 _30404_ (.A(_01677_),
    .B(_01680_),
    .Y(_01899_));
 sky130_fd_sc_hd__xnor2_2 _30405_ (.A(_01898_),
    .B(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__and3_2 _30406_ (.A(_01778_),
    .B(_01779_),
    .C(_01900_),
    .X(_01901_));
 sky130_fd_sc_hd__a21oi_2 _30407_ (.A1(_01778_),
    .A2(_01779_),
    .B1(_01900_),
    .Y(_01902_));
 sky130_fd_sc_hd__a211o_2 _30408_ (.A1(_01682_),
    .A2(_01684_),
    .B1(_01901_),
    .C1(_01902_),
    .X(_01903_));
 sky130_fd_sc_hd__o211ai_2 _30409_ (.A1(_01901_),
    .A2(_01902_),
    .B1(_01682_),
    .C1(_01684_),
    .Y(_01904_));
 sky130_fd_sc_hd__o211ai_2 _30410_ (.A1(_01553_),
    .A2(_01555_),
    .B1(_01903_),
    .C1(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__a211o_2 _30411_ (.A1(_01903_),
    .A2(_01904_),
    .B1(_01553_),
    .C1(_01555_),
    .X(_01906_));
 sky130_fd_sc_hd__o211ai_2 _30412_ (.A1(_01686_),
    .A2(_01688_),
    .B1(_01905_),
    .C1(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__a211o_2 _30413_ (.A1(_01905_),
    .A2(_01906_),
    .B1(_01686_),
    .C1(_01688_),
    .X(_01909_));
 sky130_fd_sc_hd__nand3_2 _30414_ (.A(_01691_),
    .B(_01907_),
    .C(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__a21o_2 _30415_ (.A1(_01907_),
    .A2(_01909_),
    .B1(_01691_),
    .X(_01911_));
 sky130_fd_sc_hd__nand2_4 _30416_ (.A(_01910_),
    .B(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__o21a_2 _30417_ (.A1(_00709_),
    .A2(_01122_),
    .B1(_01694_),
    .X(_01913_));
 sky130_fd_sc_hd__o21a_2 _30418_ (.A1(_01123_),
    .A2(_01132_),
    .B1(_01913_),
    .X(_01914_));
 sky130_fd_sc_hd__nor2_2 _30419_ (.A(_01693_),
    .B(_01914_),
    .Y(_01915_));
 sky130_fd_sc_hd__xor2_2 _30420_ (.A(_01912_),
    .B(_01915_),
    .X(_01916_));
 sky130_fd_sc_hd__o21ai_2 _30421_ (.A1(_01504_),
    .A2(_01297_),
    .B1(_01503_),
    .Y(_01917_));
 sky130_fd_sc_hd__and2b_2 _30422_ (.A_N(_01492_),
    .B(_01493_),
    .X(_01918_));
 sky130_fd_sc_hd__and2b_2 _30423_ (.A_N(_01495_),
    .B(_01494_),
    .X(_01920_));
 sky130_fd_sc_hd__and3_2 _30424_ (.A(_01394_),
    .B(_01395_),
    .C(_01397_),
    .X(_01921_));
 sky130_fd_sc_hd__and2b_2 _30425_ (.A_N(_01353_),
    .B(_01352_),
    .X(_01922_));
 sky130_fd_sc_hd__or2b_2 _30426_ (.A(_01383_),
    .B_N(_01391_),
    .X(_01923_));
 sky130_fd_sc_hd__and4_2 _30427_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[49]),
    .D(iX[50]),
    .X(_01924_));
 sky130_fd_sc_hd__a22oi_2 _30428_ (.A1(iY[45]),
    .A2(iX[49]),
    .B1(iX[50]),
    .B2(iY[44]),
    .Y(_01925_));
 sky130_fd_sc_hd__nor2_2 _30429_ (.A(_01924_),
    .B(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2_2 _30430_ (.A(iY[46]),
    .B(iX[48]),
    .Y(_01927_));
 sky130_fd_sc_hd__xnor2_2 _30431_ (.A(_01926_),
    .B(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__and4_2 _30432_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[52]),
    .D(iX[53]),
    .X(_01929_));
 sky130_fd_sc_hd__a22oi_2 _30433_ (.A1(iY[42]),
    .A2(iX[52]),
    .B1(iX[53]),
    .B2(iY[41]),
    .Y(_01931_));
 sky130_fd_sc_hd__nor2_2 _30434_ (.A(_01929_),
    .B(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__nand2_2 _30435_ (.A(iY[43]),
    .B(iX[51]),
    .Y(_01933_));
 sky130_fd_sc_hd__xnor2_2 _30436_ (.A(_01932_),
    .B(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__o21ba_2 _30437_ (.A1(_01349_),
    .A2(_01351_),
    .B1_N(_01347_),
    .X(_01935_));
 sky130_fd_sc_hd__xnor2_2 _30438_ (.A(_01934_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__and2_2 _30439_ (.A(_01928_),
    .B(_01936_),
    .X(_01937_));
 sky130_fd_sc_hd__nor2_2 _30440_ (.A(_01928_),
    .B(_01936_),
    .Y(_01938_));
 sky130_fd_sc_hd__or2_2 _30441_ (.A(_01937_),
    .B(_01938_),
    .X(_01939_));
 sky130_fd_sc_hd__a21o_2 _30442_ (.A1(_01389_),
    .A2(_01923_),
    .B1(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__nand3_2 _30443_ (.A(_01389_),
    .B(_01923_),
    .C(_01939_),
    .Y(_01942_));
 sky130_fd_sc_hd__o211ai_2 _30444_ (.A1(_01922_),
    .A2(_01355_),
    .B1(_01940_),
    .C1(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__a211o_2 _30445_ (.A1(_01940_),
    .A2(_01942_),
    .B1(_01922_),
    .C1(_01355_),
    .X(_01944_));
 sky130_fd_sc_hd__or2b_2 _30446_ (.A(_01371_),
    .B_N(_01369_),
    .X(_01945_));
 sky130_fd_sc_hd__nand2_2 _30447_ (.A(_01372_),
    .B(_01378_),
    .Y(_01946_));
 sky130_fd_sc_hd__and4_2 _30448_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[59]),
    .D(iX[60]),
    .X(_01947_));
 sky130_fd_sc_hd__a22oi_2 _30449_ (.A1(iY[35]),
    .A2(iX[59]),
    .B1(iX[60]),
    .B2(iY[34]),
    .Y(_01948_));
 sky130_fd_sc_hd__nor2_2 _30450_ (.A(_01947_),
    .B(_01948_),
    .Y(_01949_));
 sky130_fd_sc_hd__nand2_2 _30451_ (.A(iY[33]),
    .B(iX[61]),
    .Y(_01950_));
 sky130_fd_sc_hd__xnor2_2 _30452_ (.A(_01949_),
    .B(_01950_),
    .Y(_01951_));
 sky130_fd_sc_hd__o21ba_2 _30453_ (.A1(_01366_),
    .A2(_01368_),
    .B1_N(_01365_),
    .X(_01953_));
 sky130_fd_sc_hd__xnor2_2 _30454_ (.A(_01951_),
    .B(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__and2_2 _30455_ (.A(iY[36]),
    .B(iX[62]),
    .X(_01955_));
 sky130_fd_sc_hd__and3_2 _30456_ (.A(iY[32]),
    .B(iX[58]),
    .C(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__a22oi_2 _30457_ (.A1(iY[36]),
    .A2(iX[58]),
    .B1(iX[62]),
    .B2(iY[32]),
    .Y(_01957_));
 sky130_fd_sc_hd__o2bb2a_2 _30458_ (.A1_N(iY[37]),
    .A2_N(iX[57]),
    .B1(_01956_),
    .B2(_01957_),
    .X(_01958_));
 sky130_fd_sc_hd__and4bb_2 _30459_ (.A_N(_01956_),
    .B_N(_01957_),
    .C(iY[37]),
    .D(iX[57]),
    .X(_01959_));
 sky130_fd_sc_hd__nor2_2 _30460_ (.A(_01958_),
    .B(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__xnor2_2 _30461_ (.A(_01954_),
    .B(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__a21o_2 _30462_ (.A1(_01945_),
    .A2(_01946_),
    .B1(_01961_),
    .X(_01962_));
 sky130_fd_sc_hd__nand3_2 _30463_ (.A(_01945_),
    .B(_01946_),
    .C(_01961_),
    .Y(_01964_));
 sky130_fd_sc_hd__o21ba_2 _30464_ (.A1(_01385_),
    .A2(_01387_),
    .B1_N(_01384_),
    .X(_01965_));
 sky130_fd_sc_hd__and4_2 _30465_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[55]),
    .D(iX[56]),
    .X(_01966_));
 sky130_fd_sc_hd__a22oi_2 _30466_ (.A1(iY[39]),
    .A2(iX[55]),
    .B1(iX[56]),
    .B2(iY[38]),
    .Y(_01967_));
 sky130_fd_sc_hd__nor2_2 _30467_ (.A(_01966_),
    .B(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_2 _30468_ (.A(iY[40]),
    .B(iX[54]),
    .Y(_01969_));
 sky130_fd_sc_hd__xnor2_2 _30469_ (.A(_01968_),
    .B(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__o21ai_2 _30470_ (.A1(_01374_),
    .A2(_01377_),
    .B1(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__or3_2 _30471_ (.A(_01374_),
    .B(_01377_),
    .C(_01970_),
    .X(_01972_));
 sky130_fd_sc_hd__and2_2 _30472_ (.A(_01971_),
    .B(_01972_),
    .X(_01973_));
 sky130_fd_sc_hd__xnor2_2 _30473_ (.A(_01965_),
    .B(_01973_),
    .Y(_01975_));
 sky130_fd_sc_hd__nand3_2 _30474_ (.A(_01962_),
    .B(_01964_),
    .C(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__a21o_2 _30475_ (.A1(_01962_),
    .A2(_01964_),
    .B1(_01975_),
    .X(_01977_));
 sky130_fd_sc_hd__nand2_2 _30476_ (.A(_01380_),
    .B(_01394_),
    .Y(_01978_));
 sky130_fd_sc_hd__and3_2 _30477_ (.A(_01976_),
    .B(_01977_),
    .C(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__a21oi_2 _30478_ (.A1(_01976_),
    .A2(_01977_),
    .B1(_01978_),
    .Y(_01980_));
 sky130_fd_sc_hd__nor2_2 _30479_ (.A(_01979_),
    .B(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__a21o_2 _30480_ (.A1(_01943_),
    .A2(_01944_),
    .B1(_01981_),
    .X(_01982_));
 sky130_fd_sc_hd__and3_2 _30481_ (.A(_01981_),
    .B(_01943_),
    .C(_01944_),
    .X(_01983_));
 sky130_fd_sc_hd__inv_2 _30482_ (.A(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__o211ai_2 _30483_ (.A1(_01921_),
    .A2(_01400_),
    .B1(_01982_),
    .C1(_01984_),
    .Y(_01986_));
 sky130_fd_sc_hd__a211o_2 _30484_ (.A1(_01982_),
    .A2(_01984_),
    .B1(_01921_),
    .C1(_01400_),
    .X(_01987_));
 sky130_fd_sc_hd__nand2_2 _30485_ (.A(_01986_),
    .B(_01987_),
    .Y(_01988_));
 sky130_fd_sc_hd__inv_2 _30486_ (.A(_01437_),
    .Y(_01989_));
 sky130_fd_sc_hd__and4_2 _30487_ (.A(iX[40]),
    .B(iX[41]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_01990_));
 sky130_fd_sc_hd__a22oi_2 _30488_ (.A1(iX[41]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[40]),
    .Y(_01991_));
 sky130_fd_sc_hd__nor2_2 _30489_ (.A(_01990_),
    .B(_01991_),
    .Y(_01992_));
 sky130_fd_sc_hd__nand2_2 _30490_ (.A(iX[39]),
    .B(iY[55]),
    .Y(_01993_));
 sky130_fd_sc_hd__xnor2_2 _30491_ (.A(_01992_),
    .B(_01993_),
    .Y(_01994_));
 sky130_fd_sc_hd__and4_2 _30492_ (.A(iX[43]),
    .B(iX[44]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_01995_));
 sky130_fd_sc_hd__a22oi_2 _30493_ (.A1(iX[44]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[43]),
    .Y(_01996_));
 sky130_fd_sc_hd__nor2_2 _30494_ (.A(_01995_),
    .B(_01996_),
    .Y(_01997_));
 sky130_fd_sc_hd__nand2_2 _30495_ (.A(iX[42]),
    .B(iY[52]),
    .Y(_01998_));
 sky130_fd_sc_hd__xnor2_2 _30496_ (.A(_01997_),
    .B(_01998_),
    .Y(_01999_));
 sky130_fd_sc_hd__o21ba_2 _30497_ (.A1(_01413_),
    .A2(_01416_),
    .B1_N(_01412_),
    .X(_02000_));
 sky130_fd_sc_hd__xnor2_2 _30498_ (.A(_01999_),
    .B(_02000_),
    .Y(_02001_));
 sky130_fd_sc_hd__and2_2 _30499_ (.A(_01994_),
    .B(_02001_),
    .X(_02002_));
 sky130_fd_sc_hd__nor2_2 _30500_ (.A(_01994_),
    .B(_02001_),
    .Y(_02003_));
 sky130_fd_sc_hd__or2_2 _30501_ (.A(_02002_),
    .B(_02003_),
    .X(_02004_));
 sky130_fd_sc_hd__or3_2 _30502_ (.A(_01424_),
    .B(_01429_),
    .C(_01430_),
    .X(_02005_));
 sky130_fd_sc_hd__o21ba_2 _30503_ (.A1(_01343_),
    .A2(_01345_),
    .B1_N(_01342_),
    .X(_02007_));
 sky130_fd_sc_hd__and4_2 _30504_ (.A(iX[46]),
    .B(iX[47]),
    .C(iY[47]),
    .D(iY[48]),
    .X(_02008_));
 sky130_fd_sc_hd__a22oi_2 _30505_ (.A1(iX[47]),
    .A2(iY[47]),
    .B1(iY[48]),
    .B2(iX[46]),
    .Y(_02009_));
 sky130_fd_sc_hd__nand2_2 _30506_ (.A(iX[45]),
    .B(iY[49]),
    .Y(_02010_));
 sky130_fd_sc_hd__o21a_2 _30507_ (.A1(_02008_),
    .A2(_02009_),
    .B1(_02010_),
    .X(_02011_));
 sky130_fd_sc_hd__nor3_2 _30508_ (.A(_02008_),
    .B(_02009_),
    .C(_02010_),
    .Y(_02012_));
 sky130_fd_sc_hd__nor2_2 _30509_ (.A(_02011_),
    .B(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__xnor2_2 _30510_ (.A(_02007_),
    .B(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__o21ai_2 _30511_ (.A1(_01426_),
    .A2(_01430_),
    .B1(_02014_),
    .Y(_02015_));
 sky130_fd_sc_hd__or3_2 _30512_ (.A(_01426_),
    .B(_01430_),
    .C(_02014_),
    .X(_02016_));
 sky130_fd_sc_hd__nand2_2 _30513_ (.A(_02015_),
    .B(_02016_),
    .Y(_02018_));
 sky130_fd_sc_hd__a21oi_2 _30514_ (.A1(_02005_),
    .A2(_01433_),
    .B1(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__and3_2 _30515_ (.A(_02005_),
    .B(_01433_),
    .C(_02018_),
    .X(_02020_));
 sky130_fd_sc_hd__or3_2 _30516_ (.A(_02004_),
    .B(_02019_),
    .C(_02020_),
    .X(_02021_));
 sky130_fd_sc_hd__o21ai_2 _30517_ (.A1(_02019_),
    .A2(_02020_),
    .B1(_02004_),
    .Y(_02022_));
 sky130_fd_sc_hd__nand2_2 _30518_ (.A(_02021_),
    .B(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__a21oi_2 _30519_ (.A1(_01358_),
    .A2(_01361_),
    .B1(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__and3_2 _30520_ (.A(_01358_),
    .B(_01361_),
    .C(_02023_),
    .X(_02025_));
 sky130_fd_sc_hd__a211oi_2 _30521_ (.A1(_01989_),
    .A2(_01439_),
    .B1(_02024_),
    .C1(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__o211a_2 _30522_ (.A1(_02024_),
    .A2(_02025_),
    .B1(_01989_),
    .C1(_01439_),
    .X(_02027_));
 sky130_fd_sc_hd__or3_2 _30523_ (.A(_01988_),
    .B(_02026_),
    .C(_02027_),
    .X(_02029_));
 sky130_fd_sc_hd__inv_2 _30524_ (.A(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__o21a_2 _30525_ (.A1(_02026_),
    .A2(_02027_),
    .B1(_01988_),
    .X(_02031_));
 sky130_fd_sc_hd__a211oi_2 _30526_ (.A1(_01402_),
    .A2(_01446_),
    .B1(_02030_),
    .C1(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__o211a_2 _30527_ (.A1(_02030_),
    .A2(_02031_),
    .B1(_01402_),
    .C1(_01446_),
    .X(_02033_));
 sky130_fd_sc_hd__inv_2 _30528_ (.A(_01482_),
    .Y(_02034_));
 sky130_fd_sc_hd__and4_2 _30529_ (.A(iX[34]),
    .B(iX[35]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_02035_));
 sky130_fd_sc_hd__a22oi_2 _30530_ (.A1(iX[35]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[34]),
    .Y(_02036_));
 sky130_fd_sc_hd__nor2_2 _30531_ (.A(_02035_),
    .B(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__nand2_2 _30532_ (.A(iX[33]),
    .B(iY[61]),
    .Y(_02038_));
 sky130_fd_sc_hd__xnor2_2 _30533_ (.A(_02037_),
    .B(_02038_),
    .Y(_02040_));
 sky130_fd_sc_hd__o21ba_2 _30534_ (.A1(_01455_),
    .A2(_01457_),
    .B1_N(_01454_),
    .X(_02041_));
 sky130_fd_sc_hd__xnor2_2 _30535_ (.A(_02040_),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__nand3_2 _30536_ (.A(iX[32]),
    .B(iY[62]),
    .C(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__a21o_2 _30537_ (.A1(iX[32]),
    .A2(iY[62]),
    .B1(_02042_),
    .X(_02044_));
 sky130_fd_sc_hd__nand2_2 _30538_ (.A(_02043_),
    .B(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__nor2_2 _30539_ (.A(_01460_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__and2_2 _30540_ (.A(_01460_),
    .B(_02045_),
    .X(_02047_));
 sky130_fd_sc_hd__or2_2 _30541_ (.A(_02046_),
    .B(_02047_),
    .X(_02048_));
 sky130_fd_sc_hd__or2b_2 _30542_ (.A(_01467_),
    .B_N(_01473_),
    .X(_02049_));
 sky130_fd_sc_hd__or2b_2 _30543_ (.A(_01466_),
    .B_N(_01474_),
    .X(_02051_));
 sky130_fd_sc_hd__and2b_2 _30544_ (.A_N(_01418_),
    .B(_01417_),
    .X(_02052_));
 sky130_fd_sc_hd__o21ba_2 _30545_ (.A1(_01470_),
    .A2(_01472_),
    .B1_N(_01468_),
    .X(_02053_));
 sky130_fd_sc_hd__o21ba_2 _30546_ (.A1(_01408_),
    .A2(_01410_),
    .B1_N(_01407_),
    .X(_02054_));
 sky130_fd_sc_hd__and4_2 _30547_ (.A(iX[37]),
    .B(iX[38]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_02055_));
 sky130_fd_sc_hd__a22oi_2 _30548_ (.A1(iX[38]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[37]),
    .Y(_02056_));
 sky130_fd_sc_hd__nor2_2 _30549_ (.A(_02055_),
    .B(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__nand2_2 _30550_ (.A(iX[36]),
    .B(iY[58]),
    .Y(_02058_));
 sky130_fd_sc_hd__xnor2_2 _30551_ (.A(_02057_),
    .B(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__xnor2_2 _30552_ (.A(_02054_),
    .B(_02059_),
    .Y(_02060_));
 sky130_fd_sc_hd__xnor2_2 _30553_ (.A(_02053_),
    .B(_02060_),
    .Y(_02062_));
 sky130_fd_sc_hd__o21a_2 _30554_ (.A1(_02052_),
    .A2(_01420_),
    .B1(_02062_),
    .X(_02063_));
 sky130_fd_sc_hd__nor3_2 _30555_ (.A(_02052_),
    .B(_01420_),
    .C(_02062_),
    .Y(_02064_));
 sky130_fd_sc_hd__a211oi_2 _30556_ (.A1(_02049_),
    .A2(_02051_),
    .B1(_02063_),
    .C1(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__o211a_2 _30557_ (.A1(_02063_),
    .A2(_02064_),
    .B1(_02049_),
    .C1(_02051_),
    .X(_02066_));
 sky130_fd_sc_hd__nor2_2 _30558_ (.A(_02065_),
    .B(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__o21a_2 _30559_ (.A1(_01476_),
    .A2(_01478_),
    .B1(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__nor3_2 _30560_ (.A(_01476_),
    .B(_01478_),
    .C(_02067_),
    .Y(_02069_));
 sky130_fd_sc_hd__or3_2 _30561_ (.A(_02048_),
    .B(_02068_),
    .C(_02069_),
    .X(_02070_));
 sky130_fd_sc_hd__o21ai_2 _30562_ (.A1(_02068_),
    .A2(_02069_),
    .B1(_02048_),
    .Y(_02071_));
 sky130_fd_sc_hd__o211a_2 _30563_ (.A1(_01442_),
    .A2(_01444_),
    .B1(_02070_),
    .C1(_02071_),
    .X(_02073_));
 sky130_fd_sc_hd__a211oi_2 _30564_ (.A1(_02070_),
    .A2(_02071_),
    .B1(_01442_),
    .C1(_01444_),
    .Y(_02074_));
 sky130_fd_sc_hd__or2_2 _30565_ (.A(_02073_),
    .B(_02074_),
    .X(_02075_));
 sky130_fd_sc_hd__a21oi_2 _30566_ (.A1(_02034_),
    .A2(_01484_),
    .B1(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hd__and3_2 _30567_ (.A(_02034_),
    .B(_01484_),
    .C(_02075_),
    .X(_02077_));
 sky130_fd_sc_hd__nor4_2 _30568_ (.A(_02032_),
    .B(_02033_),
    .C(_02076_),
    .D(_02077_),
    .Y(_02078_));
 sky130_fd_sc_hd__o22a_2 _30569_ (.A1(_02032_),
    .A2(_02033_),
    .B1(_02076_),
    .B2(_02077_),
    .X(_02079_));
 sky130_fd_sc_hd__nor2_2 _30570_ (.A(_02078_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__a21o_2 _30571_ (.A1(_01453_),
    .A2(_01490_),
    .B1(_01451_),
    .X(_02081_));
 sky130_fd_sc_hd__xor2_2 _30572_ (.A(_02080_),
    .B(_02081_),
    .X(_02082_));
 sky130_fd_sc_hd__nor2_2 _30573_ (.A(_01486_),
    .B(_01488_),
    .Y(_02084_));
 sky130_fd_sc_hd__xnor2_2 _30574_ (.A(_02082_),
    .B(_02084_),
    .Y(_02085_));
 sky130_fd_sc_hd__o21ai_2 _30575_ (.A1(_01918_),
    .A2(_01920_),
    .B1(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__or3_2 _30576_ (.A(_01918_),
    .B(_01920_),
    .C(_02085_),
    .X(_02087_));
 sky130_fd_sc_hd__and3_2 _30577_ (.A(_01497_),
    .B(_02086_),
    .C(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__and2_2 _30578_ (.A(_02086_),
    .B(_02087_),
    .X(_02089_));
 sky130_fd_sc_hd__nor2_2 _30579_ (.A(_01497_),
    .B(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__or2_2 _30580_ (.A(_02088_),
    .B(_02090_),
    .X(_02091_));
 sky130_fd_sc_hd__a21oi_2 _30581_ (.A1(_01500_),
    .A2(_01917_),
    .B1(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__and3_2 _30582_ (.A(_01500_),
    .B(_01917_),
    .C(_02091_),
    .X(_02093_));
 sky130_fd_sc_hd__nor2_2 _30583_ (.A(_02092_),
    .B(_02093_),
    .Y(_02095_));
 sky130_fd_sc_hd__xor2_2 _30584_ (.A(_01916_),
    .B(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__xor2_2 _30585_ (.A(oO[30]),
    .B(_02096_),
    .X(_02097_));
 sky130_fd_sc_hd__or2b_2 _30586_ (.A(_01506_),
    .B_N(_01698_),
    .X(_02098_));
 sky130_fd_sc_hd__a21boi_2 _30587_ (.A1(_10830_),
    .A2(_01699_),
    .B1_N(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__xnor2_2 _30588_ (.A(_02097_),
    .B(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__a211o_2 _30589_ (.A1(_01706_),
    .A2(_01730_),
    .B1(_02100_),
    .C1(_01702_),
    .X(_02101_));
 sky130_fd_sc_hd__a21o_2 _30590_ (.A1(_01706_),
    .A2(_01730_),
    .B1(_01702_),
    .X(_02102_));
 sky130_fd_sc_hd__nand2_2 _30591_ (.A(_02100_),
    .B(_02102_),
    .Y(_02103_));
 sky130_fd_sc_hd__and2_2 _30592_ (.A(_02101_),
    .B(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__xor2_2 _30593_ (.A(_01729_),
    .B(_02104_),
    .X(_02106_));
 sky130_fd_sc_hd__a311o_2 _30594_ (.A1(_01308_),
    .A2(_01715_),
    .A3(_01709_),
    .B1(_01712_),
    .C1(_02106_),
    .X(_02107_));
 sky130_fd_sc_hd__a31o_2 _30595_ (.A1(_01308_),
    .A2(_01715_),
    .A3(_01709_),
    .B1(_01712_),
    .X(_02108_));
 sky130_fd_sc_hd__nand2_2 _30596_ (.A(_02106_),
    .B(_02108_),
    .Y(_02109_));
 sky130_fd_sc_hd__and2_2 _30597_ (.A(_02107_),
    .B(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__buf_1 _30598_ (.A(_02110_),
    .X(oO[62]));
 sky130_fd_sc_hd__or2_2 _30599_ (.A(_02097_),
    .B(_02099_),
    .X(_02111_));
 sky130_fd_sc_hd__or2b_2 _30600_ (.A(oO[30]),
    .B_N(_02096_),
    .X(_02112_));
 sky130_fd_sc_hd__o21ai_2 _30601_ (.A1(_01916_),
    .A2(_02095_),
    .B1(_02112_),
    .Y(_02113_));
 sky130_fd_sc_hd__and2b_2 _30602_ (.A_N(_01935_),
    .B(_01934_),
    .X(_02114_));
 sky130_fd_sc_hd__or2b_2 _30603_ (.A(_01965_),
    .B_N(_01973_),
    .X(_02116_));
 sky130_fd_sc_hd__and4_2 _30604_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[50]),
    .D(iX[51]),
    .X(_02117_));
 sky130_fd_sc_hd__a22oi_2 _30605_ (.A1(iY[45]),
    .A2(iX[50]),
    .B1(iX[51]),
    .B2(iY[44]),
    .Y(_02118_));
 sky130_fd_sc_hd__nor2_2 _30606_ (.A(_02117_),
    .B(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_2 _30607_ (.A(iY[46]),
    .B(iX[49]),
    .Y(_02120_));
 sky130_fd_sc_hd__xnor2_2 _30608_ (.A(_02119_),
    .B(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__and4_2 _30609_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[53]),
    .D(iX[54]),
    .X(_02122_));
 sky130_fd_sc_hd__a22oi_2 _30610_ (.A1(iY[42]),
    .A2(iX[53]),
    .B1(iX[54]),
    .B2(iY[41]),
    .Y(_02123_));
 sky130_fd_sc_hd__nor2_2 _30611_ (.A(_02122_),
    .B(_02123_),
    .Y(_02124_));
 sky130_fd_sc_hd__nand2_2 _30612_ (.A(iY[43]),
    .B(iX[52]),
    .Y(_02125_));
 sky130_fd_sc_hd__xnor2_2 _30613_ (.A(_02124_),
    .B(_02125_),
    .Y(_02127_));
 sky130_fd_sc_hd__o21ba_2 _30614_ (.A1(_01931_),
    .A2(_01933_),
    .B1_N(_01929_),
    .X(_02128_));
 sky130_fd_sc_hd__xnor2_2 _30615_ (.A(_02127_),
    .B(_02128_),
    .Y(_02129_));
 sky130_fd_sc_hd__and2_2 _30616_ (.A(_02121_),
    .B(_02129_),
    .X(_02130_));
 sky130_fd_sc_hd__nor2_2 _30617_ (.A(_02121_),
    .B(_02129_),
    .Y(_02131_));
 sky130_fd_sc_hd__or2_2 _30618_ (.A(_02130_),
    .B(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__a21o_2 _30619_ (.A1(_01971_),
    .A2(_02116_),
    .B1(_02132_),
    .X(_02133_));
 sky130_fd_sc_hd__nand3_2 _30620_ (.A(_01971_),
    .B(_02116_),
    .C(_02132_),
    .Y(_02134_));
 sky130_fd_sc_hd__o211ai_2 _30621_ (.A1(_02114_),
    .A2(_01937_),
    .B1(_02133_),
    .C1(_02134_),
    .Y(_02135_));
 sky130_fd_sc_hd__a211o_2 _30622_ (.A1(_02133_),
    .A2(_02134_),
    .B1(_02114_),
    .C1(_01937_),
    .X(_02136_));
 sky130_fd_sc_hd__or2b_2 _30623_ (.A(_01953_),
    .B_N(_01951_),
    .X(_02138_));
 sky130_fd_sc_hd__nand2_2 _30624_ (.A(_01954_),
    .B(_01960_),
    .Y(_02139_));
 sky130_fd_sc_hd__and4_2 _30625_ (.A(iY[34]),
    .B(iY[35]),
    .C(iX[60]),
    .D(iX[61]),
    .X(_02140_));
 sky130_fd_sc_hd__a22oi_2 _30626_ (.A1(iY[35]),
    .A2(iX[60]),
    .B1(iX[61]),
    .B2(iY[34]),
    .Y(_02141_));
 sky130_fd_sc_hd__nor2_2 _30627_ (.A(_02140_),
    .B(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__a21oi_2 _30628_ (.A1(iY[33]),
    .A2(iX[62]),
    .B1(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__and3_2 _30629_ (.A(iY[33]),
    .B(iX[62]),
    .C(_02142_),
    .X(_02144_));
 sky130_fd_sc_hd__nor2_2 _30630_ (.A(_02143_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__o21ba_2 _30631_ (.A1(_01948_),
    .A2(_01950_),
    .B1_N(_01947_),
    .X(_02146_));
 sky130_fd_sc_hd__xnor2_2 _30632_ (.A(_02145_),
    .B(_02146_),
    .Y(_02147_));
 sky130_fd_sc_hd__and3_2 _30633_ (.A(iY[32]),
    .B(iX[63]),
    .C(_00730_),
    .X(_02149_));
 sky130_fd_sc_hd__a21oi_2 _30634_ (.A1(iY[32]),
    .A2(iX[63]),
    .B1(_00730_),
    .Y(_02150_));
 sky130_fd_sc_hd__o2bb2a_2 _30635_ (.A1_N(iY[37]),
    .A2_N(iX[58]),
    .B1(_02149_),
    .B2(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__and4bb_2 _30636_ (.A_N(_02149_),
    .B_N(_02150_),
    .C(iY[37]),
    .D(iX[58]),
    .X(_02152_));
 sky130_fd_sc_hd__nor2_2 _30637_ (.A(_02151_),
    .B(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__xnor2_2 _30638_ (.A(_02147_),
    .B(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__a21o_2 _30639_ (.A1(_02138_),
    .A2(_02139_),
    .B1(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__nand3_2 _30640_ (.A(_02138_),
    .B(_02139_),
    .C(_02154_),
    .Y(_02156_));
 sky130_fd_sc_hd__o21ba_2 _30641_ (.A1(_01967_),
    .A2(_01969_),
    .B1_N(_01966_),
    .X(_02157_));
 sky130_fd_sc_hd__nand2_2 _30642_ (.A(iY[39]),
    .B(iX[56]),
    .Y(_02158_));
 sky130_fd_sc_hd__nand2_2 _30643_ (.A(iY[38]),
    .B(iX[57]),
    .Y(_02160_));
 sky130_fd_sc_hd__and4_2 _30644_ (.A(iY[38]),
    .B(iY[39]),
    .C(iX[56]),
    .D(iX[57]),
    .X(_02161_));
 sky130_fd_sc_hd__a21oi_2 _30645_ (.A1(_02158_),
    .A2(_02160_),
    .B1(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__nand2_2 _30646_ (.A(iY[40]),
    .B(iX[55]),
    .Y(_02163_));
 sky130_fd_sc_hd__xnor2_2 _30647_ (.A(_02162_),
    .B(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hd__o21ai_2 _30648_ (.A1(_01956_),
    .A2(_01959_),
    .B1(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__or3_2 _30649_ (.A(_01956_),
    .B(_01959_),
    .C(_02164_),
    .X(_02166_));
 sky130_fd_sc_hd__and2_2 _30650_ (.A(_02165_),
    .B(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__xnor2_2 _30651_ (.A(_02157_),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__nand3_2 _30652_ (.A(_02155_),
    .B(_02156_),
    .C(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__a21o_2 _30653_ (.A1(_02155_),
    .A2(_02156_),
    .B1(_02168_),
    .X(_02171_));
 sky130_fd_sc_hd__nand2_2 _30654_ (.A(_01962_),
    .B(_01976_),
    .Y(_02172_));
 sky130_fd_sc_hd__and3_2 _30655_ (.A(_02169_),
    .B(_02171_),
    .C(_02172_),
    .X(_02173_));
 sky130_fd_sc_hd__a21oi_2 _30656_ (.A1(_02169_),
    .A2(_02171_),
    .B1(_02172_),
    .Y(_02174_));
 sky130_fd_sc_hd__nor2_2 _30657_ (.A(_02173_),
    .B(_02174_),
    .Y(_02175_));
 sky130_fd_sc_hd__a21o_2 _30658_ (.A1(_02135_),
    .A2(_02136_),
    .B1(_02175_),
    .X(_02176_));
 sky130_fd_sc_hd__and3_2 _30659_ (.A(_02175_),
    .B(_02135_),
    .C(_02136_),
    .X(_02177_));
 sky130_fd_sc_hd__inv_2 _30660_ (.A(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__o211ai_2 _30661_ (.A1(_01979_),
    .A2(_01983_),
    .B1(_02176_),
    .C1(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hd__a211o_2 _30662_ (.A1(_02176_),
    .A2(_02178_),
    .B1(_01979_),
    .C1(_01983_),
    .X(_02180_));
 sky130_fd_sc_hd__nand2_2 _30663_ (.A(_02179_),
    .B(_02180_),
    .Y(_02182_));
 sky130_fd_sc_hd__inv_2 _30664_ (.A(_02019_),
    .Y(_02183_));
 sky130_fd_sc_hd__and4_2 _30665_ (.A(iX[41]),
    .B(iX[42]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_02184_));
 sky130_fd_sc_hd__a22oi_2 _30666_ (.A1(iX[42]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[41]),
    .Y(_02185_));
 sky130_fd_sc_hd__nor2_2 _30667_ (.A(_02184_),
    .B(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__nand2_2 _30668_ (.A(iX[40]),
    .B(iY[55]),
    .Y(_02187_));
 sky130_fd_sc_hd__xnor2_2 _30669_ (.A(_02186_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__and4_2 _30670_ (.A(iX[44]),
    .B(iX[45]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_02189_));
 sky130_fd_sc_hd__a22oi_2 _30671_ (.A1(iX[45]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[44]),
    .Y(_02190_));
 sky130_fd_sc_hd__nor2_2 _30672_ (.A(_02189_),
    .B(_02190_),
    .Y(_02191_));
 sky130_fd_sc_hd__nand2_2 _30673_ (.A(iX[43]),
    .B(iY[52]),
    .Y(_02193_));
 sky130_fd_sc_hd__xnor2_2 _30674_ (.A(_02191_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__o21ba_2 _30675_ (.A1(_01996_),
    .A2(_01998_),
    .B1_N(_01995_),
    .X(_02195_));
 sky130_fd_sc_hd__xnor2_2 _30676_ (.A(_02194_),
    .B(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__and2_2 _30677_ (.A(_02188_),
    .B(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__nor2_2 _30678_ (.A(_02188_),
    .B(_02196_),
    .Y(_02198_));
 sky130_fd_sc_hd__or2_2 _30679_ (.A(_02197_),
    .B(_02198_),
    .X(_02199_));
 sky130_fd_sc_hd__or3_2 _30680_ (.A(_02007_),
    .B(_02011_),
    .C(_02012_),
    .X(_02200_));
 sky130_fd_sc_hd__o21ba_2 _30681_ (.A1(_01925_),
    .A2(_01927_),
    .B1_N(_01924_),
    .X(_02201_));
 sky130_fd_sc_hd__and4_2 _30682_ (.A(iX[47]),
    .B(iY[47]),
    .C(iX[48]),
    .D(iY[48]),
    .X(_02202_));
 sky130_fd_sc_hd__a22oi_2 _30683_ (.A1(iY[47]),
    .A2(iX[48]),
    .B1(iY[48]),
    .B2(iX[47]),
    .Y(_02204_));
 sky130_fd_sc_hd__nand2_2 _30684_ (.A(iX[46]),
    .B(iY[49]),
    .Y(_02205_));
 sky130_fd_sc_hd__o21a_2 _30685_ (.A1(_02202_),
    .A2(_02204_),
    .B1(_02205_),
    .X(_02206_));
 sky130_fd_sc_hd__nor3_2 _30686_ (.A(_02202_),
    .B(_02204_),
    .C(_02205_),
    .Y(_02207_));
 sky130_fd_sc_hd__nor2_2 _30687_ (.A(_02206_),
    .B(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__xnor2_2 _30688_ (.A(_02201_),
    .B(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__o21ai_2 _30689_ (.A1(_02008_),
    .A2(_02012_),
    .B1(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__or3_2 _30690_ (.A(_02008_),
    .B(_02012_),
    .C(_02209_),
    .X(_02211_));
 sky130_fd_sc_hd__nand2_2 _30691_ (.A(_02210_),
    .B(_02211_),
    .Y(_02212_));
 sky130_fd_sc_hd__a21oi_2 _30692_ (.A1(_02200_),
    .A2(_02015_),
    .B1(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__and3_2 _30693_ (.A(_02200_),
    .B(_02015_),
    .C(_02212_),
    .X(_02215_));
 sky130_fd_sc_hd__or3_2 _30694_ (.A(_02199_),
    .B(_02213_),
    .C(_02215_),
    .X(_02216_));
 sky130_fd_sc_hd__o21ai_2 _30695_ (.A1(_02213_),
    .A2(_02215_),
    .B1(_02199_),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_2 _30696_ (.A(_02216_),
    .B(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__a21oi_2 _30697_ (.A1(_01940_),
    .A2(_01943_),
    .B1(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__and3_2 _30698_ (.A(_01940_),
    .B(_01943_),
    .C(_02218_),
    .X(_02220_));
 sky130_fd_sc_hd__a211oi_2 _30699_ (.A1(_02183_),
    .A2(_02021_),
    .B1(_02219_),
    .C1(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__o211a_2 _30700_ (.A1(_02219_),
    .A2(_02220_),
    .B1(_02183_),
    .C1(_02021_),
    .X(_02222_));
 sky130_fd_sc_hd__or3_2 _30701_ (.A(_02182_),
    .B(_02221_),
    .C(_02222_),
    .X(_02223_));
 sky130_fd_sc_hd__inv_2 _30702_ (.A(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__o21a_2 _30703_ (.A1(_02221_),
    .A2(_02222_),
    .B1(_02182_),
    .X(_02226_));
 sky130_fd_sc_hd__a211oi_2 _30704_ (.A1(_01986_),
    .A2(_02029_),
    .B1(_02224_),
    .C1(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__o211a_2 _30705_ (.A1(_02224_),
    .A2(_02226_),
    .B1(_01986_),
    .C1(_02029_),
    .X(_02228_));
 sky130_fd_sc_hd__or2_2 _30706_ (.A(_02227_),
    .B(_02228_),
    .X(_02229_));
 sky130_fd_sc_hd__inv_2 _30707_ (.A(_02068_),
    .Y(_02230_));
 sky130_fd_sc_hd__or2b_2 _30708_ (.A(_02041_),
    .B_N(_02040_),
    .X(_02231_));
 sky130_fd_sc_hd__and4_2 _30709_ (.A(iX[35]),
    .B(iX[36]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_02232_));
 sky130_fd_sc_hd__a22oi_2 _30710_ (.A1(iX[36]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[35]),
    .Y(_02233_));
 sky130_fd_sc_hd__nor2_2 _30711_ (.A(_02232_),
    .B(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__nand2_2 _30712_ (.A(iX[34]),
    .B(iY[61]),
    .Y(_02235_));
 sky130_fd_sc_hd__xnor2_2 _30713_ (.A(_02234_),
    .B(_02235_),
    .Y(_02237_));
 sky130_fd_sc_hd__o21ba_2 _30714_ (.A1(_02036_),
    .A2(_02038_),
    .B1_N(_02035_),
    .X(_02238_));
 sky130_fd_sc_hd__xnor2_2 _30715_ (.A(_02237_),
    .B(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__and2_2 _30716_ (.A(iX[33]),
    .B(iY[62]),
    .X(_02240_));
 sky130_fd_sc_hd__or2_2 _30717_ (.A(_02239_),
    .B(_02240_),
    .X(_02241_));
 sky130_fd_sc_hd__nand2_2 _30718_ (.A(_02239_),
    .B(_02240_),
    .Y(_02242_));
 sky130_fd_sc_hd__nand2_2 _30719_ (.A(_02241_),
    .B(_02242_),
    .Y(_02243_));
 sky130_fd_sc_hd__a21oi_2 _30720_ (.A1(_02231_),
    .A2(_02043_),
    .B1(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__and3_2 _30721_ (.A(_02231_),
    .B(_02043_),
    .C(_02243_),
    .X(_02245_));
 sky130_fd_sc_hd__nor2_2 _30722_ (.A(_02244_),
    .B(_02245_),
    .Y(_02246_));
 sky130_fd_sc_hd__nand2_2 _30723_ (.A(iX[32]),
    .B(iY[63]),
    .Y(_02248_));
 sky130_fd_sc_hd__xnor2_2 _30724_ (.A(_02246_),
    .B(_02248_),
    .Y(_02249_));
 sky130_fd_sc_hd__or2b_2 _30725_ (.A(_02054_),
    .B_N(_02059_),
    .X(_02250_));
 sky130_fd_sc_hd__or2b_2 _30726_ (.A(_02053_),
    .B_N(_02060_),
    .X(_02251_));
 sky130_fd_sc_hd__and2b_2 _30727_ (.A_N(_02000_),
    .B(_01999_),
    .X(_02252_));
 sky130_fd_sc_hd__o21ba_2 _30728_ (.A1(_02056_),
    .A2(_02058_),
    .B1_N(_02055_),
    .X(_02253_));
 sky130_fd_sc_hd__o21ba_2 _30729_ (.A1(_01991_),
    .A2(_01993_),
    .B1_N(_01990_),
    .X(_02254_));
 sky130_fd_sc_hd__and4_2 _30730_ (.A(iX[38]),
    .B(iX[39]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_02255_));
 sky130_fd_sc_hd__a22oi_2 _30731_ (.A1(iX[39]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[38]),
    .Y(_02256_));
 sky130_fd_sc_hd__nor2_2 _30732_ (.A(_02255_),
    .B(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__nand2_2 _30733_ (.A(iX[37]),
    .B(iY[58]),
    .Y(_02259_));
 sky130_fd_sc_hd__xnor2_2 _30734_ (.A(_02257_),
    .B(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hd__xnor2_2 _30735_ (.A(_02254_),
    .B(_02260_),
    .Y(_02261_));
 sky130_fd_sc_hd__xnor2_2 _30736_ (.A(_02253_),
    .B(_02261_),
    .Y(_02262_));
 sky130_fd_sc_hd__o21a_2 _30737_ (.A1(_02252_),
    .A2(_02002_),
    .B1(_02262_),
    .X(_02263_));
 sky130_fd_sc_hd__nor3_2 _30738_ (.A(_02252_),
    .B(_02002_),
    .C(_02262_),
    .Y(_02264_));
 sky130_fd_sc_hd__a211oi_2 _30739_ (.A1(_02250_),
    .A2(_02251_),
    .B1(_02263_),
    .C1(_02264_),
    .Y(_02265_));
 sky130_fd_sc_hd__o211a_2 _30740_ (.A1(_02263_),
    .A2(_02264_),
    .B1(_02250_),
    .C1(_02251_),
    .X(_02266_));
 sky130_fd_sc_hd__nor2_2 _30741_ (.A(_02063_),
    .B(_02065_),
    .Y(_02267_));
 sky130_fd_sc_hd__or3_2 _30742_ (.A(_02265_),
    .B(_02266_),
    .C(_02267_),
    .X(_02268_));
 sky130_fd_sc_hd__o21ai_2 _30743_ (.A1(_02265_),
    .A2(_02266_),
    .B1(_02267_),
    .Y(_02270_));
 sky130_fd_sc_hd__and3_2 _30744_ (.A(_02249_),
    .B(_02268_),
    .C(_02270_),
    .X(_02271_));
 sky130_fd_sc_hd__a21oi_2 _30745_ (.A1(_02268_),
    .A2(_02270_),
    .B1(_02249_),
    .Y(_02272_));
 sky130_fd_sc_hd__nor2_2 _30746_ (.A(_02271_),
    .B(_02272_),
    .Y(_02273_));
 sky130_fd_sc_hd__o21a_2 _30747_ (.A1(_02024_),
    .A2(_02026_),
    .B1(_02273_),
    .X(_02274_));
 sky130_fd_sc_hd__nor3_2 _30748_ (.A(_02024_),
    .B(_02026_),
    .C(_02273_),
    .Y(_02275_));
 sky130_fd_sc_hd__a211oi_2 _30749_ (.A1(_02230_),
    .A2(_02070_),
    .B1(_02274_),
    .C1(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__o211a_2 _30750_ (.A1(_02274_),
    .A2(_02275_),
    .B1(_02230_),
    .C1(_02070_),
    .X(_02277_));
 sky130_fd_sc_hd__nor2_2 _30751_ (.A(_02276_),
    .B(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__xnor2_2 _30752_ (.A(_02229_),
    .B(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__o21ai_2 _30753_ (.A1(_02032_),
    .A2(_02078_),
    .B1(_02279_),
    .Y(_02281_));
 sky130_fd_sc_hd__or3_2 _30754_ (.A(_02032_),
    .B(_02078_),
    .C(_02279_),
    .X(_02282_));
 sky130_fd_sc_hd__o211ai_2 _30755_ (.A1(_02073_),
    .A2(_02076_),
    .B1(_02281_),
    .C1(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__a211o_2 _30756_ (.A1(_02281_),
    .A2(_02282_),
    .B1(_02073_),
    .C1(_02076_),
    .X(_02284_));
 sky130_fd_sc_hd__and2b_2 _30757_ (.A_N(_02084_),
    .B(_02082_),
    .X(_02285_));
 sky130_fd_sc_hd__a21o_2 _30758_ (.A1(_02080_),
    .A2(_02081_),
    .B1(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__and3_2 _30759_ (.A(_02283_),
    .B(_02284_),
    .C(_02286_),
    .X(_02287_));
 sky130_fd_sc_hd__a21o_2 _30760_ (.A1(_02283_),
    .A2(_02284_),
    .B1(_02286_),
    .X(_02288_));
 sky130_fd_sc_hd__and2b_2 _30761_ (.A_N(_02287_),
    .B(_02288_),
    .X(_02289_));
 sky130_fd_sc_hd__xor2_2 _30762_ (.A(_02046_),
    .B(_02289_),
    .X(_02290_));
 sky130_fd_sc_hd__xnor2_2 _30763_ (.A(_02086_),
    .B(_02290_),
    .Y(_02292_));
 sky130_fd_sc_hd__or2_2 _30764_ (.A(_02088_),
    .B(_02092_),
    .X(_02293_));
 sky130_fd_sc_hd__xnor2_2 _30765_ (.A(_02292_),
    .B(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__o31a_2 _30766_ (.A1(_01693_),
    .A2(_01912_),
    .A3(_01914_),
    .B1(_01910_),
    .X(_02295_));
 sky130_fd_sc_hd__and2b_2 _30767_ (.A_N(_01526_),
    .B(_01748_),
    .X(_02296_));
 sky130_fd_sc_hd__nand2_2 _30768_ (.A(_01775_),
    .B(_01778_),
    .Y(_02297_));
 sky130_fd_sc_hd__xnor2_2 _30769_ (.A(_02296_),
    .B(_02297_),
    .Y(_02298_));
 sky130_fd_sc_hd__and2b_2 _30770_ (.A_N(_01899_),
    .B(_01898_),
    .X(_02299_));
 sky130_fd_sc_hd__nand2_2 _30771_ (.A(_01771_),
    .B(_01773_),
    .Y(_02300_));
 sky130_fd_sc_hd__and2b_2 _30772_ (.A_N(_01822_),
    .B(_01783_),
    .X(_02301_));
 sky130_fd_sc_hd__and2b_2 _30773_ (.A_N(_01823_),
    .B(_01781_),
    .X(_02303_));
 sky130_fd_sc_hd__nor2_2 _30774_ (.A(_01737_),
    .B(_01738_),
    .Y(_02304_));
 sky130_fd_sc_hd__and2b_2 _30775_ (.A_N(_01739_),
    .B(_01747_),
    .X(_02305_));
 sky130_fd_sc_hd__or4_4 _30776_ (.A(_18120_),
    .B(_16271_),
    .C(_01512_),
    .D(_00943_),
    .X(_02306_));
 sky130_fd_sc_hd__a22o_2 _30777_ (.A1(_14629_),
    .A2(_00565_),
    .B1(_01510_),
    .B2(_18749_),
    .X(_02307_));
 sky130_fd_sc_hd__and4_2 _30778_ (.A(_15616_),
    .B(_01521_),
    .C(_02306_),
    .D(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__a22oi_2 _30779_ (.A1(_15616_),
    .A2(_01521_),
    .B1(_02306_),
    .B2(_02307_),
    .Y(_02309_));
 sky130_fd_sc_hd__or2_2 _30780_ (.A(_02308_),
    .B(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__buf_1 _30781_ (.A(_01512_),
    .X(_02311_));
 sky130_fd_sc_hd__or3_2 _30782_ (.A(_18120_),
    .B(_02311_),
    .C(_01511_),
    .X(_02312_));
 sky130_fd_sc_hd__o21a_2 _30783_ (.A1(_01734_),
    .A2(_01736_),
    .B1(_02312_),
    .X(_02314_));
 sky130_fd_sc_hd__xnor2_2 _30784_ (.A(_02310_),
    .B(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__buf_1 _30785_ (.A(_01746_),
    .X(_02316_));
 sky130_fd_sc_hd__buf_1 _30786_ (.A(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__nand2_2 _30787_ (.A(iY[31]),
    .B(iY[63]),
    .Y(_02318_));
 sky130_fd_sc_hd__or2_2 _30788_ (.A(iY[31]),
    .B(iY[63]),
    .X(_02319_));
 sky130_fd_sc_hd__nand2_2 _30789_ (.A(_02318_),
    .B(_02319_),
    .Y(_02320_));
 sky130_fd_sc_hd__a21boi_2 _30790_ (.A1(_01741_),
    .A2(_01745_),
    .B1_N(_01740_),
    .Y(_02321_));
 sky130_fd_sc_hd__xnor2_2 _30791_ (.A(_02320_),
    .B(_02321_),
    .Y(_02322_));
 sky130_fd_sc_hd__o22a_2 _30792_ (.A1(_11571_),
    .A2(_02317_),
    .B1(_02322_),
    .B2(_11579_),
    .X(_02323_));
 sky130_fd_sc_hd__or3b_2 _30793_ (.A(_11571_),
    .B(_02322_),
    .C_N(_01747_),
    .X(_02325_));
 sky130_fd_sc_hd__or2b_2 _30794_ (.A(_02323_),
    .B_N(_02325_),
    .X(_02326_));
 sky130_fd_sc_hd__xor2_2 _30795_ (.A(_02315_),
    .B(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__o21ai_2 _30796_ (.A1(_02304_),
    .A2(_02305_),
    .B1(_02327_),
    .Y(_02328_));
 sky130_fd_sc_hd__or3_2 _30797_ (.A(_02304_),
    .B(_02305_),
    .C(_02327_),
    .X(_02329_));
 sky130_fd_sc_hd__nand3_2 _30798_ (.A(_01751_),
    .B(_01767_),
    .C(_01768_),
    .Y(_02330_));
 sky130_fd_sc_hd__nand2_2 _30799_ (.A(_01762_),
    .B(_01764_),
    .Y(_02331_));
 sky130_fd_sc_hd__nor2_2 _30800_ (.A(_01800_),
    .B(_01801_),
    .Y(_02332_));
 sky130_fd_sc_hd__a21o_2 _30801_ (.A1(_01792_),
    .A2(_01802_),
    .B1(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__nand2_2 _30802_ (.A(_01758_),
    .B(_01761_),
    .Y(_02334_));
 sky130_fd_sc_hd__o21bai_2 _30803_ (.A1(_01788_),
    .A2(_01789_),
    .B1_N(_01786_),
    .Y(_02336_));
 sky130_fd_sc_hd__or4b_2 _30804_ (.A(_00195_),
    .B(_00589_),
    .C(_18343_),
    .D_N(_18729_),
    .X(_02337_));
 sky130_fd_sc_hd__buf_1 _30805_ (.A(_16277_),
    .X(_02338_));
 sky130_fd_sc_hd__a22o_2 _30806_ (.A1(_02338_),
    .A2(_18734_),
    .B1(_18729_),
    .B2(_01564_),
    .X(_02339_));
 sky130_fd_sc_hd__a22o_2 _30807_ (.A1(_18754_),
    .A2(_01757_),
    .B1(_02337_),
    .B2(_02339_),
    .X(_02340_));
 sky130_fd_sc_hd__nand4_2 _30808_ (.A(_18754_),
    .B(_01757_),
    .C(_02337_),
    .D(_02339_),
    .Y(_02341_));
 sky130_fd_sc_hd__nand3_2 _30809_ (.A(_02336_),
    .B(_02340_),
    .C(_02341_),
    .Y(_02342_));
 sky130_fd_sc_hd__a21o_2 _30810_ (.A1(_02340_),
    .A2(_02341_),
    .B1(_02336_),
    .X(_02343_));
 sky130_fd_sc_hd__nand3_2 _30811_ (.A(_02334_),
    .B(_02342_),
    .C(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__a21o_2 _30812_ (.A1(_02342_),
    .A2(_02343_),
    .B1(_02334_),
    .X(_02345_));
 sky130_fd_sc_hd__nand3_2 _30813_ (.A(_02333_),
    .B(_02344_),
    .C(_02345_),
    .Y(_02347_));
 sky130_fd_sc_hd__a21o_2 _30814_ (.A1(_02344_),
    .A2(_02345_),
    .B1(_02333_),
    .X(_02348_));
 sky130_fd_sc_hd__and3_2 _30815_ (.A(_02331_),
    .B(_02347_),
    .C(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__a21oi_2 _30816_ (.A1(_02347_),
    .A2(_02348_),
    .B1(_02331_),
    .Y(_02350_));
 sky130_fd_sc_hd__a211o_2 _30817_ (.A1(_01767_),
    .A2(_02330_),
    .B1(_02349_),
    .C1(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__o211ai_2 _30818_ (.A1(_02349_),
    .A2(_02350_),
    .B1(_01767_),
    .C1(_02330_),
    .Y(_02352_));
 sky130_fd_sc_hd__nand4_2 _30819_ (.A(_02328_),
    .B(_02329_),
    .C(_02351_),
    .D(_02352_),
    .Y(_02353_));
 sky130_fd_sc_hd__a22o_2 _30820_ (.A1(_02328_),
    .A2(_02329_),
    .B1(_02351_),
    .B2(_02352_),
    .X(_02354_));
 sky130_fd_sc_hd__o211ai_2 _30821_ (.A1(_02301_),
    .A2(_02303_),
    .B1(_02353_),
    .C1(_02354_),
    .Y(_02355_));
 sky130_fd_sc_hd__a211o_2 _30822_ (.A1(_02353_),
    .A2(_02354_),
    .B1(_02301_),
    .C1(_02303_),
    .X(_02356_));
 sky130_fd_sc_hd__nand3_2 _30823_ (.A(_02300_),
    .B(_02355_),
    .C(_02356_),
    .Y(_02358_));
 sky130_fd_sc_hd__a21o_2 _30824_ (.A1(_02355_),
    .A2(_02356_),
    .B1(_02300_),
    .X(_02359_));
 sky130_fd_sc_hd__or2_2 _30825_ (.A(_01894_),
    .B(_01895_),
    .X(_02360_));
 sky130_fd_sc_hd__or2_2 _30826_ (.A(_01824_),
    .B(_01896_),
    .X(_02361_));
 sky130_fd_sc_hd__nor2_2 _30827_ (.A(_01891_),
    .B(_01892_),
    .Y(_02362_));
 sky130_fd_sc_hd__and2_2 _30828_ (.A(_01848_),
    .B(_01893_),
    .X(_02363_));
 sky130_fd_sc_hd__o21ai_2 _30829_ (.A1(_01834_),
    .A2(_01845_),
    .B1(_01843_),
    .Y(_02364_));
 sky130_fd_sc_hd__and2_2 _30830_ (.A(_01850_),
    .B(_01857_),
    .X(_02365_));
 sky130_fd_sc_hd__nand2_2 _30831_ (.A(_14605_),
    .B(_17488_),
    .Y(_02366_));
 sky130_fd_sc_hd__or3_2 _30832_ (.A(_01605_),
    .B(_00255_),
    .C(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__a22o_2 _30833_ (.A1(_14606_),
    .A2(_17006_),
    .B1(_17488_),
    .B2(_14411_),
    .X(_02369_));
 sky130_fd_sc_hd__nand2_2 _30834_ (.A(_02367_),
    .B(_02369_),
    .Y(_02370_));
 sky130_fd_sc_hd__nor2_2 _30835_ (.A(_15173_),
    .B(_01828_),
    .Y(_02371_));
 sky130_fd_sc_hd__xor2_2 _30836_ (.A(_02370_),
    .B(_02371_),
    .X(_02372_));
 sky130_fd_sc_hd__nor2_2 _30837_ (.A(_13893_),
    .B(_17482_),
    .Y(_02373_));
 sky130_fd_sc_hd__nor2_2 _30838_ (.A(_18791_),
    .B(_18443_),
    .Y(_02374_));
 sky130_fd_sc_hd__xnor2_2 _30839_ (.A(_02373_),
    .B(_02374_),
    .Y(_02375_));
 sky130_fd_sc_hd__nand2_2 _30840_ (.A(_01039_),
    .B(_17702_),
    .Y(_02376_));
 sky130_fd_sc_hd__xnor2_2 _30841_ (.A(_02375_),
    .B(_02376_),
    .Y(_02377_));
 sky130_fd_sc_hd__nand2_2 _30842_ (.A(_01611_),
    .B(_01835_),
    .Y(_02378_));
 sky130_fd_sc_hd__o21a_2 _30843_ (.A1(_01836_),
    .A2(_01838_),
    .B1(_02378_),
    .X(_02380_));
 sky130_fd_sc_hd__xnor2_2 _30844_ (.A(_02377_),
    .B(_02380_),
    .Y(_02381_));
 sky130_fd_sc_hd__xor2_2 _30845_ (.A(_02372_),
    .B(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__o21ai_2 _30846_ (.A1(_02365_),
    .A2(_01859_),
    .B1(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__or3_2 _30847_ (.A(_02365_),
    .B(_01859_),
    .C(_02382_),
    .X(_02384_));
 sky130_fd_sc_hd__nand2_2 _30848_ (.A(_02383_),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__xnor2_2 _30849_ (.A(_02364_),
    .B(_02385_),
    .Y(_02386_));
 sky130_fd_sc_hd__or2_2 _30850_ (.A(_01888_),
    .B(_01889_),
    .X(_02387_));
 sky130_fd_sc_hd__or2_2 _30851_ (.A(_01861_),
    .B(_01890_),
    .X(_02388_));
 sky130_fd_sc_hd__or2_2 _30852_ (.A(_01655_),
    .B(_01657_),
    .X(_02389_));
 sky130_fd_sc_hd__buf_1 _30853_ (.A(_02389_),
    .X(_02391_));
 sky130_fd_sc_hd__nor2_2 _30854_ (.A(_11794_),
    .B(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__nand3_2 _30855_ (.A(_11585_),
    .B(_01880_),
    .C(_01881_),
    .Y(_02393_));
 sky130_fd_sc_hd__nand2_2 _30856_ (.A(iX[31]),
    .B(iX[63]),
    .Y(_02394_));
 sky130_fd_sc_hd__or2_2 _30857_ (.A(iX[31]),
    .B(iX[63]),
    .X(_02395_));
 sky130_fd_sc_hd__nand2_2 _30858_ (.A(_02394_),
    .B(_02395_),
    .Y(_02396_));
 sky130_fd_sc_hd__and3_2 _30859_ (.A(_01877_),
    .B(_01880_),
    .C(_02396_),
    .X(_02397_));
 sky130_fd_sc_hd__a21oi_2 _30860_ (.A1(_01877_),
    .A2(_01880_),
    .B1(_02396_),
    .Y(_02398_));
 sky130_fd_sc_hd__or4_4 _30861_ (.A(_11567_),
    .B(_02393_),
    .C(_02397_),
    .D(_02398_),
    .X(_02399_));
 sky130_fd_sc_hd__o31ai_2 _30862_ (.A1(_11567_),
    .A2(_02397_),
    .A3(_02398_),
    .B1(_02393_),
    .Y(_02400_));
 sky130_fd_sc_hd__nand3_2 _30863_ (.A(_02392_),
    .B(_02399_),
    .C(_02400_),
    .Y(_02402_));
 sky130_fd_sc_hd__a21o_2 _30864_ (.A1(_02399_),
    .A2(_02400_),
    .B1(_02392_),
    .X(_02403_));
 sky130_fd_sc_hd__or3_2 _30865_ (.A(_11567_),
    .B(_02389_),
    .C(_02393_),
    .X(_02404_));
 sky130_fd_sc_hd__a21bo_2 _30866_ (.A1(_01871_),
    .A2(_01883_),
    .B1_N(_02404_),
    .X(_02405_));
 sky130_fd_sc_hd__and3_2 _30867_ (.A(_02402_),
    .B(_02403_),
    .C(_02405_),
    .X(_02406_));
 sky130_fd_sc_hd__a21oi_2 _30868_ (.A1(_02402_),
    .A2(_02403_),
    .B1(_02405_),
    .Y(_02407_));
 sky130_fd_sc_hd__nand2_2 _30869_ (.A(_15887_),
    .B(_01643_),
    .Y(_02408_));
 sky130_fd_sc_hd__nor2_2 _30870_ (.A(_15650_),
    .B(_01087_),
    .Y(_02409_));
 sky130_fd_sc_hd__and3_2 _30871_ (.A(_00661_),
    .B(_01650_),
    .C(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__a21oi_2 _30872_ (.A1(_00661_),
    .A2(_01650_),
    .B1(_02409_),
    .Y(_02411_));
 sky130_fd_sc_hd__nor2_2 _30873_ (.A(_02410_),
    .B(_02411_),
    .Y(_02413_));
 sky130_fd_sc_hd__xnor2_2 _30874_ (.A(_02408_),
    .B(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__or3b_2 _30875_ (.A(_02406_),
    .B(_02407_),
    .C_N(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__o21bai_2 _30876_ (.A1(_02406_),
    .A2(_02407_),
    .B1_N(_02414_),
    .Y(_02416_));
 sky130_fd_sc_hd__nor2_2 _30877_ (.A(_01884_),
    .B(_01885_),
    .Y(_02417_));
 sky130_fd_sc_hd__a21o_2 _30878_ (.A1(_01870_),
    .A2(_01887_),
    .B1(_02417_),
    .X(_02418_));
 sky130_fd_sc_hd__and3_2 _30879_ (.A(_02415_),
    .B(_02416_),
    .C(_02418_),
    .X(_02419_));
 sky130_fd_sc_hd__a21oi_2 _30880_ (.A1(_02415_),
    .A2(_02416_),
    .B1(_02418_),
    .Y(_02420_));
 sky130_fd_sc_hd__or2b_2 _30881_ (.A(_01851_),
    .B_N(_01856_),
    .X(_02421_));
 sky130_fd_sc_hd__a31o_2 _30882_ (.A1(_18192_),
    .A2(_01862_),
    .A3(_01868_),
    .B1(_01867_),
    .X(_02422_));
 sky130_fd_sc_hd__o22a_2 _30883_ (.A1(_12852_),
    .A2(_00271_),
    .B1(_00666_),
    .B2(_12848_),
    .X(_02424_));
 sky130_fd_sc_hd__a31o_2 _30884_ (.A1(_14637_),
    .A2(_01862_),
    .A3(_01852_),
    .B1(_02424_),
    .X(_02425_));
 sky130_fd_sc_hd__nor2_2 _30885_ (.A(_14626_),
    .B(_01066_),
    .Y(_02426_));
 sky130_fd_sc_hd__xnor2_2 _30886_ (.A(_02425_),
    .B(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__xnor2_2 _30887_ (.A(_02422_),
    .B(_02427_),
    .Y(_02428_));
 sky130_fd_sc_hd__a21oi_2 _30888_ (.A1(_01854_),
    .A2(_02421_),
    .B1(_02428_),
    .Y(_02429_));
 sky130_fd_sc_hd__and3_2 _30889_ (.A(_01854_),
    .B(_02421_),
    .C(_02428_),
    .X(_02430_));
 sky130_fd_sc_hd__nor2_2 _30890_ (.A(_02429_),
    .B(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__nor3b_2 _30891_ (.A(_02419_),
    .B(_02420_),
    .C_N(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__o21ba_2 _30892_ (.A1(_02419_),
    .A2(_02420_),
    .B1_N(_02431_),
    .X(_02433_));
 sky130_fd_sc_hd__a211o_2 _30893_ (.A1(_02387_),
    .A2(_02388_),
    .B1(_02432_),
    .C1(_02433_),
    .X(_02435_));
 sky130_fd_sc_hd__o211ai_2 _30894_ (.A1(_02432_),
    .A2(_02433_),
    .B1(_02387_),
    .C1(_02388_),
    .Y(_02436_));
 sky130_fd_sc_hd__nand3_2 _30895_ (.A(_02386_),
    .B(_02435_),
    .C(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__a21o_2 _30896_ (.A1(_02435_),
    .A2(_02436_),
    .B1(_02386_),
    .X(_02438_));
 sky130_fd_sc_hd__o211a_2 _30897_ (.A1(_02362_),
    .A2(_02363_),
    .B1(_02437_),
    .C1(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__a211oi_2 _30898_ (.A1(_02437_),
    .A2(_02438_),
    .B1(_02362_),
    .C1(_02363_),
    .Y(_02440_));
 sky130_fd_sc_hd__and2b_2 _30899_ (.A_N(_01819_),
    .B(_01816_),
    .X(_02441_));
 sky130_fd_sc_hd__a21o_2 _30900_ (.A1(_01803_),
    .A2(_01821_),
    .B1(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__or2b_2 _30901_ (.A(_01847_),
    .B_N(_01825_),
    .X(_02443_));
 sky130_fd_sc_hd__a21bo_2 _30902_ (.A1(_01826_),
    .A2(_01846_),
    .B1_N(_02443_),
    .X(_02444_));
 sky130_fd_sc_hd__and4_2 _30903_ (.A(_01785_),
    .B(_00999_),
    .C(_17630_),
    .D(_18101_),
    .X(_02446_));
 sky130_fd_sc_hd__o22a_2 _30904_ (.A1(_01797_),
    .A2(_17408_),
    .B1(_17627_),
    .B2(_16288_),
    .X(_02447_));
 sky130_fd_sc_hd__nor2_2 _30905_ (.A(_02446_),
    .B(_02447_),
    .Y(_02448_));
 sky130_fd_sc_hd__nand2_2 _30906_ (.A(_01784_),
    .B(_18326_),
    .Y(_02449_));
 sky130_fd_sc_hd__xor2_2 _30907_ (.A(_02448_),
    .B(_02449_),
    .X(_02450_));
 sky130_fd_sc_hd__or3b_2 _30908_ (.A(_15005_),
    .B(_16617_),
    .C_N(_01793_),
    .X(_02451_));
 sky130_fd_sc_hd__a2bb2o_2 _30909_ (.A1_N(_15005_),
    .A2_N(_16257_),
    .B1(_16613_),
    .B2(_15888_),
    .X(_02452_));
 sky130_fd_sc_hd__nand2_2 _30910_ (.A(_02451_),
    .B(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__or2_2 _30911_ (.A(_15648_),
    .B(_18363_),
    .X(_02454_));
 sky130_fd_sc_hd__xnor2_2 _30912_ (.A(_02453_),
    .B(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__o21a_2 _30913_ (.A1(_01796_),
    .A2(_01799_),
    .B1(_01794_),
    .X(_02457_));
 sky130_fd_sc_hd__xnor2_2 _30914_ (.A(_02455_),
    .B(_02457_),
    .Y(_02458_));
 sky130_fd_sc_hd__or2_2 _30915_ (.A(_02450_),
    .B(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__nand2_2 _30916_ (.A(_02450_),
    .B(_02458_),
    .Y(_02460_));
 sky130_fd_sc_hd__and2_2 _30917_ (.A(_02459_),
    .B(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__or2_2 _30918_ (.A(_00996_),
    .B(_01810_),
    .X(_02462_));
 sky130_fd_sc_hd__buf_1 _30919_ (.A(_15005_),
    .X(_02463_));
 sky130_fd_sc_hd__o22a_2 _30920_ (.A1(_01807_),
    .A2(_01808_),
    .B1(_02462_),
    .B2(_02463_),
    .X(_02464_));
 sky130_fd_sc_hd__a21oi_2 _30921_ (.A1(_01830_),
    .A2(_01833_),
    .B1(_01827_),
    .Y(_02465_));
 sky130_fd_sc_hd__or2_2 _30922_ (.A(_15597_),
    .B(_16312_),
    .X(_02466_));
 sky130_fd_sc_hd__buf_1 _30923_ (.A(_02466_),
    .X(_02468_));
 sky130_fd_sc_hd__o22a_2 _30924_ (.A1(_18181_),
    .A2(_15598_),
    .B1(_16312_),
    .B2(_15154_),
    .X(_02469_));
 sky130_fd_sc_hd__o21ba_2 _30925_ (.A1(_01808_),
    .A2(_02468_),
    .B1_N(_02469_),
    .X(_02470_));
 sky130_fd_sc_hd__buf_1 _30926_ (.A(_14998_),
    .X(_02471_));
 sky130_fd_sc_hd__nor2_2 _30927_ (.A(_02471_),
    .B(_15835_),
    .Y(_02472_));
 sky130_fd_sc_hd__xor2_2 _30928_ (.A(_02470_),
    .B(_02472_),
    .X(_02473_));
 sky130_fd_sc_hd__xnor2_2 _30929_ (.A(_02465_),
    .B(_02473_),
    .Y(_02474_));
 sky130_fd_sc_hd__xnor2_2 _30930_ (.A(_02464_),
    .B(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__a21oi_2 _30931_ (.A1(_01806_),
    .A2(_01815_),
    .B1(_01813_),
    .Y(_02476_));
 sky130_fd_sc_hd__xnor2_2 _30932_ (.A(_02475_),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__xnor2_2 _30933_ (.A(_02461_),
    .B(_02477_),
    .Y(_02479_));
 sky130_fd_sc_hd__xnor2_2 _30934_ (.A(_02444_),
    .B(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__xor2_2 _30935_ (.A(_02442_),
    .B(_02480_),
    .X(_02481_));
 sky130_fd_sc_hd__nor3b_2 _30936_ (.A(_02439_),
    .B(_02440_),
    .C_N(_02481_),
    .Y(_02482_));
 sky130_fd_sc_hd__o21ba_2 _30937_ (.A1(_02439_),
    .A2(_02440_),
    .B1_N(_02481_),
    .X(_02483_));
 sky130_fd_sc_hd__a211o_2 _30938_ (.A1(_02360_),
    .A2(_02361_),
    .B1(_02482_),
    .C1(_02483_),
    .X(_02484_));
 sky130_fd_sc_hd__o211ai_2 _30939_ (.A1(_02482_),
    .A2(_02483_),
    .B1(_02360_),
    .C1(_02361_),
    .Y(_02485_));
 sky130_fd_sc_hd__nand4_2 _30940_ (.A(_02358_),
    .B(_02359_),
    .C(_02484_),
    .D(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__a22o_2 _30941_ (.A1(_02358_),
    .A2(_02359_),
    .B1(_02484_),
    .B2(_02485_),
    .X(_02487_));
 sky130_fd_sc_hd__o211a_2 _30942_ (.A1(_02299_),
    .A2(_01901_),
    .B1(_02486_),
    .C1(_02487_),
    .X(_02488_));
 sky130_fd_sc_hd__a211oi_2 _30943_ (.A1(_02486_),
    .A2(_02487_),
    .B1(_02299_),
    .C1(_01901_),
    .Y(_02490_));
 sky130_fd_sc_hd__nor3_2 _30944_ (.A(_02298_),
    .B(_02488_),
    .C(_02490_),
    .Y(_02491_));
 sky130_fd_sc_hd__o21a_2 _30945_ (.A1(_02488_),
    .A2(_02490_),
    .B1(_02298_),
    .X(_02492_));
 sky130_fd_sc_hd__a211o_2 _30946_ (.A1(_01903_),
    .A2(_01905_),
    .B1(_02491_),
    .C1(_02492_),
    .X(_02493_));
 sky130_fd_sc_hd__o211ai_2 _30947_ (.A1(_02491_),
    .A2(_02492_),
    .B1(_01903_),
    .C1(_01905_),
    .Y(_02494_));
 sky130_fd_sc_hd__a21boi_2 _30948_ (.A1(_02493_),
    .A2(_02494_),
    .B1_N(_01907_),
    .Y(_02495_));
 sky130_fd_sc_hd__nand3b_2 _30949_ (.A_N(_01907_),
    .B(_02493_),
    .C(_02494_),
    .Y(_02496_));
 sky130_fd_sc_hd__or2b_2 _30950_ (.A(_02495_),
    .B_N(_02496_),
    .X(_02497_));
 sky130_fd_sc_hd__xnor2_2 _30951_ (.A(_02295_),
    .B(_02497_),
    .Y(_02498_));
 sky130_fd_sc_hd__xnor2_2 _30952_ (.A(_02294_),
    .B(_02498_),
    .Y(_02499_));
 sky130_fd_sc_hd__xnor2_2 _30953_ (.A(oO[31]),
    .B(_02499_),
    .Y(_02501_));
 sky130_fd_sc_hd__xnor2_2 _30954_ (.A(_02113_),
    .B(_02501_),
    .Y(_02502_));
 sky130_fd_sc_hd__a21oi_2 _30955_ (.A1(_02111_),
    .A2(_02101_),
    .B1(_02502_),
    .Y(_02503_));
 sky130_fd_sc_hd__and3_2 _30956_ (.A(_02111_),
    .B(_02101_),
    .C(_02502_),
    .X(_02504_));
 sky130_fd_sc_hd__or2_2 _30957_ (.A(_02503_),
    .B(_02504_),
    .X(_02505_));
 sky130_fd_sc_hd__o211a_2 _30958_ (.A1(_01719_),
    .A2(_01720_),
    .B1(_01723_),
    .C1(_01727_),
    .X(_02506_));
 sky130_fd_sc_hd__nor2_2 _30959_ (.A(_02505_),
    .B(_02506_),
    .Y(_02507_));
 sky130_fd_sc_hd__nand2_2 _30960_ (.A(_02505_),
    .B(_02506_),
    .Y(_02508_));
 sky130_fd_sc_hd__and2b_2 _30961_ (.A_N(_02507_),
    .B(_02508_),
    .X(_02509_));
 sky130_fd_sc_hd__or2b_2 _30962_ (.A(_01729_),
    .B_N(_02104_),
    .X(_02510_));
 sky130_fd_sc_hd__nand2_2 _30963_ (.A(_02510_),
    .B(_02107_),
    .Y(_02512_));
 sky130_fd_sc_hd__xor2_2 _30964_ (.A(_02509_),
    .B(_02512_),
    .X(oO[63]));
 sky130_fd_sc_hd__and2_2 _30965_ (.A(_02296_),
    .B(_02297_),
    .X(_02513_));
 sky130_fd_sc_hd__a21oi_2 _30966_ (.A1(_02355_),
    .A2(_02358_),
    .B1(_02328_),
    .Y(_02514_));
 sky130_fd_sc_hd__and3_2 _30967_ (.A(_02328_),
    .B(_02355_),
    .C(_02358_),
    .X(_02515_));
 sky130_fd_sc_hd__nor2_2 _30968_ (.A(_02514_),
    .B(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__nand2_2 _30969_ (.A(_02351_),
    .B(_02353_),
    .Y(_02517_));
 sky130_fd_sc_hd__and2b_2 _30970_ (.A_N(_02479_),
    .B(_02444_),
    .X(_02518_));
 sky130_fd_sc_hd__a21o_2 _30971_ (.A1(_02442_),
    .A2(_02480_),
    .B1(_02518_),
    .X(_02519_));
 sky130_fd_sc_hd__nand2_2 _30972_ (.A(_14629_),
    .B(_01510_),
    .Y(_02520_));
 sky130_fd_sc_hd__and4_2 _30973_ (.A(_18754_),
    .B(_16268_),
    .C(_00161_),
    .D(_00565_),
    .X(_02522_));
 sky130_fd_sc_hd__a22o_2 _30974_ (.A1(_01564_),
    .A2(_00162_),
    .B1(_00565_),
    .B2(_18754_),
    .X(_02523_));
 sky130_fd_sc_hd__and2b_2 _30975_ (.A_N(_02522_),
    .B(_02523_),
    .X(_02524_));
 sky130_fd_sc_hd__xnor2_2 _30976_ (.A(_02520_),
    .B(_02524_),
    .Y(_02525_));
 sky130_fd_sc_hd__and4_2 _30977_ (.A(_18749_),
    .B(_14629_),
    .C(_00566_),
    .D(_01510_),
    .X(_02526_));
 sky130_fd_sc_hd__nor2_2 _30978_ (.A(_02526_),
    .B(_02308_),
    .Y(_02527_));
 sky130_fd_sc_hd__xnor2_2 _30979_ (.A(_02525_),
    .B(_02527_),
    .Y(_02528_));
 sky130_fd_sc_hd__nor2_2 _30980_ (.A(_11571_),
    .B(_02322_),
    .Y(_02529_));
 sky130_fd_sc_hd__nand2_2 _30981_ (.A(_18749_),
    .B(_01521_),
    .Y(_02530_));
 sky130_fd_sc_hd__nor2_2 _30982_ (.A(_16625_),
    .B(_02316_),
    .Y(_02531_));
 sky130_fd_sc_hd__xnor2_2 _30983_ (.A(_02530_),
    .B(_02531_),
    .Y(_02533_));
 sky130_fd_sc_hd__xor2_2 _30984_ (.A(_02529_),
    .B(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__xnor2_2 _30985_ (.A(_02528_),
    .B(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__o22a_2 _30986_ (.A1(_02310_),
    .A2(_02314_),
    .B1(_02315_),
    .B2(_02326_),
    .X(_02536_));
 sky130_fd_sc_hd__xor2_2 _30987_ (.A(_02535_),
    .B(_02536_),
    .X(_02537_));
 sky130_fd_sc_hd__xnor2_2 _30988_ (.A(_02325_),
    .B(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__nand2_2 _30989_ (.A(_02342_),
    .B(_02344_),
    .Y(_02539_));
 sky130_fd_sc_hd__o21ai_2 _30990_ (.A1(_02455_),
    .A2(_02457_),
    .B1(_02459_),
    .Y(_02540_));
 sky130_fd_sc_hd__nand2_2 _30991_ (.A(_02337_),
    .B(_02341_),
    .Y(_02541_));
 sky130_fd_sc_hd__o21ba_2 _30992_ (.A1(_02447_),
    .A2(_02449_),
    .B1_N(_02446_),
    .X(_02542_));
 sky130_fd_sc_hd__nand2_2 _30993_ (.A(_02338_),
    .B(_18729_),
    .Y(_02544_));
 sky130_fd_sc_hd__or3_2 _30994_ (.A(_14983_),
    .B(_18110_),
    .C(_18112_),
    .X(_02545_));
 sky130_fd_sc_hd__nand2_2 _30995_ (.A(_14652_),
    .B(_18732_),
    .Y(_02546_));
 sky130_fd_sc_hd__xor2_2 _30996_ (.A(_02545_),
    .B(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__xnor2_2 _30997_ (.A(_02544_),
    .B(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__xnor2_2 _30998_ (.A(_02542_),
    .B(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__xor2_2 _30999_ (.A(_02541_),
    .B(_02549_),
    .X(_02550_));
 sky130_fd_sc_hd__xor2_2 _31000_ (.A(_02540_),
    .B(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__xnor2_2 _31001_ (.A(_02539_),
    .B(_02551_),
    .Y(_02552_));
 sky130_fd_sc_hd__a21boi_2 _31002_ (.A1(_02331_),
    .A2(_02348_),
    .B1_N(_02347_),
    .Y(_02553_));
 sky130_fd_sc_hd__xnor2_2 _31003_ (.A(_02552_),
    .B(_02553_),
    .Y(_02555_));
 sky130_fd_sc_hd__xnor2_2 _31004_ (.A(_02538_),
    .B(_02555_),
    .Y(_02556_));
 sky130_fd_sc_hd__xnor2_2 _31005_ (.A(_02519_),
    .B(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__xnor2_2 _31006_ (.A(_02517_),
    .B(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__and2b_2 _31007_ (.A_N(_02476_),
    .B(_02475_),
    .X(_02559_));
 sky130_fd_sc_hd__a21oi_2 _31008_ (.A1(_02461_),
    .A2(_02477_),
    .B1(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__or2b_2 _31009_ (.A(_02385_),
    .B_N(_02364_),
    .X(_02561_));
 sky130_fd_sc_hd__nor2_2 _31010_ (.A(_01797_),
    .B(_17628_),
    .Y(_02562_));
 sky130_fd_sc_hd__or2_2 _31011_ (.A(_14988_),
    .B(_16922_),
    .X(_02563_));
 sky130_fd_sc_hd__or3_2 _31012_ (.A(_15648_),
    .B(_17408_),
    .C(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__o21ai_2 _31013_ (.A1(_15648_),
    .A2(_17408_),
    .B1(_02563_),
    .Y(_02566_));
 sky130_fd_sc_hd__and2_2 _31014_ (.A(_02564_),
    .B(_02566_),
    .X(_02567_));
 sky130_fd_sc_hd__xor2_2 _31015_ (.A(_02562_),
    .B(_02567_),
    .X(_02568_));
 sky130_fd_sc_hd__nor2_2 _31016_ (.A(_15005_),
    .B(_16619_),
    .Y(_02569_));
 sky130_fd_sc_hd__nor2_2 _31017_ (.A(_02471_),
    .B(_16257_),
    .Y(_02570_));
 sky130_fd_sc_hd__and3_2 _31018_ (.A(_17460_),
    .B(_16934_),
    .C(_02570_),
    .X(_02571_));
 sky130_fd_sc_hd__a21oi_2 _31019_ (.A1(_17460_),
    .A2(_16934_),
    .B1(_02570_),
    .Y(_02572_));
 sky130_fd_sc_hd__nor2_2 _31020_ (.A(_02571_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__xnor2_2 _31021_ (.A(_02569_),
    .B(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__o21a_2 _31022_ (.A1(_02453_),
    .A2(_02454_),
    .B1(_02451_),
    .X(_02575_));
 sky130_fd_sc_hd__nor2_2 _31023_ (.A(_02574_),
    .B(_02575_),
    .Y(_02577_));
 sky130_fd_sc_hd__nand2_2 _31024_ (.A(_02574_),
    .B(_02575_),
    .Y(_02578_));
 sky130_fd_sc_hd__and2b_2 _31025_ (.A_N(_02577_),
    .B(_02578_),
    .X(_02579_));
 sky130_fd_sc_hd__xnor2_2 _31026_ (.A(_02568_),
    .B(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hd__a2bb2o_2 _31027_ (.A1_N(_01808_),
    .A2_N(_02468_),
    .B1(_02470_),
    .B2(_02472_),
    .X(_02581_));
 sky130_fd_sc_hd__a21bo_2 _31028_ (.A1(_02369_),
    .A2(_02371_),
    .B1_N(_02367_),
    .X(_02582_));
 sky130_fd_sc_hd__nand2_2 _31029_ (.A(_15617_),
    .B(_16682_),
    .Y(_02583_));
 sky130_fd_sc_hd__or3_2 _31030_ (.A(_15153_),
    .B(_17696_),
    .C(_02583_),
    .X(_02584_));
 sky130_fd_sc_hd__o21ai_2 _31031_ (.A1(_16237_),
    .A2(_17696_),
    .B1(_02583_),
    .Y(_02585_));
 sky130_fd_sc_hd__and2_2 _31032_ (.A(_02584_),
    .B(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__xnor2_2 _31033_ (.A(_02468_),
    .B(_02586_),
    .Y(_02588_));
 sky130_fd_sc_hd__and2_2 _31034_ (.A(_02582_),
    .B(_02588_),
    .X(_02589_));
 sky130_fd_sc_hd__nor2_2 _31035_ (.A(_02582_),
    .B(_02588_),
    .Y(_02590_));
 sky130_fd_sc_hd__nor2_2 _31036_ (.A(_02589_),
    .B(_02590_),
    .Y(_02591_));
 sky130_fd_sc_hd__xnor2_2 _31037_ (.A(_02581_),
    .B(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__and2b_2 _31038_ (.A_N(_02473_),
    .B(_02465_),
    .X(_02593_));
 sky130_fd_sc_hd__or2b_2 _31039_ (.A(_02465_),
    .B_N(_02473_),
    .X(_02594_));
 sky130_fd_sc_hd__o21a_2 _31040_ (.A1(_02464_),
    .A2(_02593_),
    .B1(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__xnor2_2 _31041_ (.A(_02592_),
    .B(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__xnor2_2 _31042_ (.A(_02580_),
    .B(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__a21oi_2 _31043_ (.A1(_02383_),
    .A2(_02561_),
    .B1(_02597_),
    .Y(_02599_));
 sky130_fd_sc_hd__and3_2 _31044_ (.A(_02383_),
    .B(_02561_),
    .C(_02597_),
    .X(_02600_));
 sky130_fd_sc_hd__or3_2 _31045_ (.A(_02560_),
    .B(_02599_),
    .C(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__o21ai_2 _31046_ (.A1(_02599_),
    .A2(_02600_),
    .B1(_02560_),
    .Y(_02602_));
 sky130_fd_sc_hd__and2_2 _31047_ (.A(_02601_),
    .B(_02602_),
    .X(_02603_));
 sky130_fd_sc_hd__or2_2 _31048_ (.A(_02377_),
    .B(_02380_),
    .X(_02604_));
 sky130_fd_sc_hd__o21a_2 _31049_ (.A1(_02372_),
    .A2(_02381_),
    .B1(_02604_),
    .X(_02605_));
 sky130_fd_sc_hd__a21o_2 _31050_ (.A1(_02422_),
    .A2(_02427_),
    .B1(_02429_),
    .X(_02606_));
 sky130_fd_sc_hd__and4_2 _31051_ (.A(_14392_),
    .B(_14411_),
    .C(_17702_),
    .D(_18209_),
    .X(_02607_));
 sky130_fd_sc_hd__buf_1 _31052_ (.A(_13972_),
    .X(_02608_));
 sky130_fd_sc_hd__o22a_2 _31053_ (.A1(_15168_),
    .A2(_01058_),
    .B1(_18200_),
    .B2(_02608_),
    .X(_02610_));
 sky130_fd_sc_hd__nor2_2 _31054_ (.A(_02607_),
    .B(_02610_),
    .Y(_02611_));
 sky130_fd_sc_hd__xnor2_2 _31055_ (.A(_02366_),
    .B(_02611_),
    .Y(_02612_));
 sky130_fd_sc_hd__buf_1 _31056_ (.A(_13893_),
    .X(_02613_));
 sky130_fd_sc_hd__or4_2 _31057_ (.A(_14641_),
    .B(_14612_),
    .C(_18211_),
    .D(_00271_),
    .X(_02614_));
 sky130_fd_sc_hd__a22o_2 _31058_ (.A1(_13543_),
    .A2(_00662_),
    .B1(_18460_),
    .B2(_17463_),
    .X(_02615_));
 sky130_fd_sc_hd__and2_2 _31059_ (.A(_02614_),
    .B(_02615_),
    .X(_02616_));
 sky130_fd_sc_hd__or3b_2 _31060_ (.A(_02613_),
    .B(_18443_),
    .C_N(_02616_),
    .X(_02617_));
 sky130_fd_sc_hd__a21o_2 _31061_ (.A1(_13889_),
    .A2(_18463_),
    .B1(_02616_),
    .X(_02618_));
 sky130_fd_sc_hd__nand2_2 _31062_ (.A(_02617_),
    .B(_02618_),
    .Y(_02619_));
 sky130_fd_sc_hd__o2bb2ai_2 _31063_ (.A1_N(_02373_),
    .A2_N(_02374_),
    .B1(_02375_),
    .B2(_02376_),
    .Y(_02621_));
 sky130_fd_sc_hd__xnor2_2 _31064_ (.A(_02619_),
    .B(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__xnor2_2 _31065_ (.A(_02612_),
    .B(_02622_),
    .Y(_02623_));
 sky130_fd_sc_hd__xnor2_2 _31066_ (.A(_02606_),
    .B(_02623_),
    .Y(_02624_));
 sky130_fd_sc_hd__xnor2_2 _31067_ (.A(_02605_),
    .B(_02624_),
    .Y(_02625_));
 sky130_fd_sc_hd__buf_1 _31068_ (.A(_14637_),
    .X(_02626_));
 sky130_fd_sc_hd__and2b_2 _31069_ (.A_N(_02425_),
    .B(_02426_),
    .X(_02627_));
 sky130_fd_sc_hd__a31o_2 _31070_ (.A1(_02626_),
    .A2(_01862_),
    .A3(_01852_),
    .B1(_02627_),
    .X(_02628_));
 sky130_fd_sc_hd__buf_1 _31071_ (.A(_01643_),
    .X(_02629_));
 sky130_fd_sc_hd__and3_2 _31072_ (.A(_18192_),
    .B(_02629_),
    .C(_02413_),
    .X(_02630_));
 sky130_fd_sc_hd__nand2_2 _31073_ (.A(_14637_),
    .B(_01862_),
    .Y(_02632_));
 sky130_fd_sc_hd__nor3_2 _31074_ (.A(_12848_),
    .B(_01866_),
    .C(_02408_),
    .Y(_02633_));
 sky130_fd_sc_hd__a22o_2 _31075_ (.A1(_14636_),
    .A2(_01643_),
    .B1(_01650_),
    .B2(_15887_),
    .X(_02634_));
 sky130_fd_sc_hd__and2b_2 _31076_ (.A_N(_02633_),
    .B(_02634_),
    .X(_02635_));
 sky130_fd_sc_hd__xnor2_2 _31077_ (.A(_02632_),
    .B(_02635_),
    .Y(_02636_));
 sky130_fd_sc_hd__o21a_2 _31078_ (.A1(_02410_),
    .A2(_02630_),
    .B1(_02636_),
    .X(_02637_));
 sky130_fd_sc_hd__or3_2 _31079_ (.A(_02410_),
    .B(_02630_),
    .C(_02636_),
    .X(_02638_));
 sky130_fd_sc_hd__or2b_2 _31080_ (.A(_02637_),
    .B_N(_02638_),
    .X(_02639_));
 sky130_fd_sc_hd__xor2_2 _31081_ (.A(_02628_),
    .B(_02639_),
    .X(_02640_));
 sky130_fd_sc_hd__nor2_2 _31082_ (.A(_01655_),
    .B(_01657_),
    .Y(_02641_));
 sky130_fd_sc_hd__nand2_2 _31083_ (.A(_01880_),
    .B(_01881_),
    .Y(_02643_));
 sky130_fd_sc_hd__nor2_2 _31084_ (.A(_15650_),
    .B(_02643_),
    .Y(_02644_));
 sky130_fd_sc_hd__and3_2 _31085_ (.A(_15677_),
    .B(_02641_),
    .C(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__o22a_2 _31086_ (.A1(_15650_),
    .A2(_02391_),
    .B1(_02643_),
    .B2(_11794_),
    .X(_02646_));
 sky130_fd_sc_hd__buf_1 _31087_ (.A(_01087_),
    .X(_02647_));
 sky130_fd_sc_hd__inv_2 _31088_ (.A(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__and4bb_2 _31089_ (.A_N(_02645_),
    .B_N(_02646_),
    .C(_00661_),
    .D(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__o22a_2 _31090_ (.A1(_14978_),
    .A2(_02647_),
    .B1(_02645_),
    .B2(_02646_),
    .X(_02650_));
 sky130_fd_sc_hd__or2_2 _31091_ (.A(_02649_),
    .B(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__or2_2 _31092_ (.A(_02397_),
    .B(_02398_),
    .X(_02652_));
 sky130_fd_sc_hd__nor2_2 _31093_ (.A(_11576_),
    .B(_02652_),
    .Y(_02654_));
 sky130_fd_sc_hd__inv_2 _31094_ (.A(_01744_),
    .Y(_02655_));
 sky130_fd_sc_hd__o32a_2 _31095_ (.A1(_00939_),
    .A2(_00933_),
    .A3(_01519_),
    .B1(_02655_),
    .B2(_01518_),
    .X(_02656_));
 sky130_fd_sc_hd__a21bo_2 _31096_ (.A1(_01740_),
    .A2(_02318_),
    .B1_N(_02319_),
    .X(_02657_));
 sky130_fd_sc_hd__o31a_2 _31097_ (.A1(_01742_),
    .A2(_02320_),
    .A3(_02656_),
    .B1(_02657_),
    .X(_02658_));
 sky130_fd_sc_hd__or4_2 _31098_ (.A(_00939_),
    .B(_01519_),
    .C(_01742_),
    .D(_02320_),
    .X(_02659_));
 sky130_fd_sc_hd__a211o_2 _31099_ (.A1(_18336_),
    .A2(_00934_),
    .B1(_00935_),
    .C1(_02659_),
    .X(_02660_));
 sky130_fd_sc_hd__a21o_2 _31100_ (.A1(_02658_),
    .A2(_02660_),
    .B1(_11578_),
    .X(_02661_));
 sky130_fd_sc_hd__nor2_2 _31101_ (.A(iX[31]),
    .B(iX[63]),
    .Y(_02662_));
 sky130_fd_sc_hd__a31o_2 _31102_ (.A1(_01877_),
    .A2(_01880_),
    .A3(_02394_),
    .B1(_02662_),
    .X(_02663_));
 sky130_fd_sc_hd__nor2_2 _31103_ (.A(_11567_),
    .B(_02663_),
    .Y(_02665_));
 sky130_fd_sc_hd__xnor2_2 _31104_ (.A(_02661_),
    .B(_02665_),
    .Y(_02666_));
 sky130_fd_sc_hd__xor2_2 _31105_ (.A(_02654_),
    .B(_02666_),
    .X(_02667_));
 sky130_fd_sc_hd__and2_2 _31106_ (.A(_02399_),
    .B(_02402_),
    .X(_02668_));
 sky130_fd_sc_hd__xnor2_2 _31107_ (.A(_02667_),
    .B(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__xnor2_2 _31108_ (.A(_02651_),
    .B(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__nand2b_2 _31109_ (.A_N(_02406_),
    .B(_02415_),
    .Y(_02671_));
 sky130_fd_sc_hd__xor2_2 _31110_ (.A(_02670_),
    .B(_02671_),
    .X(_02672_));
 sky130_fd_sc_hd__xnor2_2 _31111_ (.A(_02640_),
    .B(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__nor2_2 _31112_ (.A(_02419_),
    .B(_02432_),
    .Y(_02674_));
 sky130_fd_sc_hd__xnor2_2 _31113_ (.A(_02673_),
    .B(_02674_),
    .Y(_02676_));
 sky130_fd_sc_hd__xnor2_2 _31114_ (.A(_02625_),
    .B(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__nand2_2 _31115_ (.A(_02435_),
    .B(_02437_),
    .Y(_02678_));
 sky130_fd_sc_hd__xnor2_2 _31116_ (.A(_02677_),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__xor2_2 _31117_ (.A(_02603_),
    .B(_02679_),
    .X(_02680_));
 sky130_fd_sc_hd__nor2_2 _31118_ (.A(_02439_),
    .B(_02482_),
    .Y(_02681_));
 sky130_fd_sc_hd__xnor2_2 _31119_ (.A(_02680_),
    .B(_02681_),
    .Y(_02682_));
 sky130_fd_sc_hd__xnor2_2 _31120_ (.A(_02558_),
    .B(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__nand2_2 _31121_ (.A(_02484_),
    .B(_02486_),
    .Y(_02684_));
 sky130_fd_sc_hd__xnor2_2 _31122_ (.A(_02683_),
    .B(_02684_),
    .Y(_02685_));
 sky130_fd_sc_hd__xor2_2 _31123_ (.A(_02516_),
    .B(_02685_),
    .X(_02687_));
 sky130_fd_sc_hd__nor2_2 _31124_ (.A(_02488_),
    .B(_02491_),
    .Y(_02688_));
 sky130_fd_sc_hd__xnor2_2 _31125_ (.A(_02687_),
    .B(_02688_),
    .Y(_02689_));
 sky130_fd_sc_hd__xor2_2 _31126_ (.A(_02513_),
    .B(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__xnor2_2 _31127_ (.A(_02493_),
    .B(_02690_),
    .Y(_02691_));
 sky130_fd_sc_hd__o21a_2 _31128_ (.A1(_01910_),
    .A2(_02495_),
    .B1(_02496_),
    .X(_02692_));
 sky130_fd_sc_hd__o41a_2 _31129_ (.A1(_01693_),
    .A2(_01912_),
    .A3(_01913_),
    .A4(_02497_),
    .B1(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__or4_4 _31130_ (.A(_01123_),
    .B(_01695_),
    .C(_01912_),
    .D(_02497_),
    .X(_02694_));
 sky130_fd_sc_hd__a21o_2 _31131_ (.A1(_01126_),
    .A2(_01131_),
    .B1(_02694_),
    .X(_02695_));
 sky130_fd_sc_hd__nand2_2 _31132_ (.A(_02693_),
    .B(_02695_),
    .Y(_02696_));
 sky130_fd_sc_hd__xnor2_2 _31133_ (.A(_02691_),
    .B(_02696_),
    .Y(_02698_));
 sky130_fd_sc_hd__or2b_2 _31134_ (.A(_02086_),
    .B_N(_02290_),
    .X(_02699_));
 sky130_fd_sc_hd__o21ai_2 _31135_ (.A1(_02088_),
    .A2(_02092_),
    .B1(_02292_),
    .Y(_02700_));
 sky130_fd_sc_hd__o21ba_2 _31136_ (.A1(_02245_),
    .A2(_02248_),
    .B1_N(_02244_),
    .X(_02701_));
 sky130_fd_sc_hd__and2b_2 _31137_ (.A_N(_02146_),
    .B(_02145_),
    .X(_02702_));
 sky130_fd_sc_hd__and2_2 _31138_ (.A(_02147_),
    .B(_02153_),
    .X(_02703_));
 sky130_fd_sc_hd__and2_2 _31139_ (.A(iY[34]),
    .B(iX[62]),
    .X(_02704_));
 sky130_fd_sc_hd__and3_2 _31140_ (.A(iY[35]),
    .B(iX[61]),
    .C(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__a21o_2 _31141_ (.A1(iY[35]),
    .A2(iX[61]),
    .B1(_02704_),
    .X(_02706_));
 sky130_fd_sc_hd__and2b_2 _31142_ (.A_N(_02705_),
    .B(_02706_),
    .X(_02707_));
 sky130_fd_sc_hd__nand2_2 _31143_ (.A(iY[33]),
    .B(iX[63]),
    .Y(_02709_));
 sky130_fd_sc_hd__xnor2_2 _31144_ (.A(_02707_),
    .B(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__nor2_2 _31145_ (.A(_02140_),
    .B(_02144_),
    .Y(_02711_));
 sky130_fd_sc_hd__xor2_2 _31146_ (.A(_02710_),
    .B(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__a22oi_2 _31147_ (.A1(iY[37]),
    .A2(iX[59]),
    .B1(iX[60]),
    .B2(iY[36]),
    .Y(_02713_));
 sky130_fd_sc_hd__and3_2 _31148_ (.A(iY[37]),
    .B(iX[60]),
    .C(_00730_),
    .X(_02714_));
 sky130_fd_sc_hd__or2_2 _31149_ (.A(_02713_),
    .B(_02714_),
    .X(_02715_));
 sky130_fd_sc_hd__xor2_2 _31150_ (.A(_02712_),
    .B(_02715_),
    .X(_02716_));
 sky130_fd_sc_hd__o21a_2 _31151_ (.A1(_02702_),
    .A2(_02703_),
    .B1(_02716_),
    .X(_02717_));
 sky130_fd_sc_hd__nor3_2 _31152_ (.A(_02702_),
    .B(_02703_),
    .C(_02716_),
    .Y(_02718_));
 sky130_fd_sc_hd__a31o_2 _31153_ (.A1(iY[40]),
    .A2(iX[55]),
    .A3(_02162_),
    .B1(_02161_),
    .X(_02720_));
 sky130_fd_sc_hd__nand2_2 _31154_ (.A(iY[39]),
    .B(iX[57]),
    .Y(_02721_));
 sky130_fd_sc_hd__nand2_2 _31155_ (.A(iY[38]),
    .B(iX[58]),
    .Y(_02722_));
 sky130_fd_sc_hd__nand2_2 _31156_ (.A(iY[39]),
    .B(iX[58]),
    .Y(_02723_));
 sky130_fd_sc_hd__nor2_2 _31157_ (.A(_02160_),
    .B(_02723_),
    .Y(_02724_));
 sky130_fd_sc_hd__a21oi_2 _31158_ (.A1(_02721_),
    .A2(_02722_),
    .B1(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__nand2_2 _31159_ (.A(iY[40]),
    .B(iX[56]),
    .Y(_02726_));
 sky130_fd_sc_hd__xnor2_2 _31160_ (.A(_02725_),
    .B(_02726_),
    .Y(_02727_));
 sky130_fd_sc_hd__o21ai_2 _31161_ (.A1(_02149_),
    .A2(_02152_),
    .B1(_02727_),
    .Y(_02728_));
 sky130_fd_sc_hd__or3_2 _31162_ (.A(_02149_),
    .B(_02152_),
    .C(_02727_),
    .X(_02729_));
 sky130_fd_sc_hd__and2_2 _31163_ (.A(_02728_),
    .B(_02729_),
    .X(_02731_));
 sky130_fd_sc_hd__xnor2_2 _31164_ (.A(_02720_),
    .B(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__nor3_2 _31165_ (.A(_02717_),
    .B(_02718_),
    .C(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hd__o21a_2 _31166_ (.A1(_02717_),
    .A2(_02718_),
    .B1(_02732_),
    .X(_02734_));
 sky130_fd_sc_hd__a211oi_2 _31167_ (.A1(_02155_),
    .A2(_02169_),
    .B1(_02733_),
    .C1(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__o211a_2 _31168_ (.A1(_02733_),
    .A2(_02734_),
    .B1(_02155_),
    .C1(_02169_),
    .X(_02736_));
 sky130_fd_sc_hd__and2b_2 _31169_ (.A_N(_02128_),
    .B(_02127_),
    .X(_02737_));
 sky130_fd_sc_hd__or2b_2 _31170_ (.A(_02157_),
    .B_N(_02167_),
    .X(_02738_));
 sky130_fd_sc_hd__and4_2 _31171_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[51]),
    .D(iX[52]),
    .X(_02739_));
 sky130_fd_sc_hd__a22oi_2 _31172_ (.A1(iY[45]),
    .A2(iX[51]),
    .B1(iX[52]),
    .B2(iY[44]),
    .Y(_02740_));
 sky130_fd_sc_hd__nor2_2 _31173_ (.A(_02739_),
    .B(_02740_),
    .Y(_02742_));
 sky130_fd_sc_hd__nand2_2 _31174_ (.A(iY[46]),
    .B(iX[50]),
    .Y(_02743_));
 sky130_fd_sc_hd__xnor2_2 _31175_ (.A(_02742_),
    .B(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hd__and4_2 _31176_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[54]),
    .D(iX[55]),
    .X(_02745_));
 sky130_fd_sc_hd__a22oi_2 _31177_ (.A1(iY[42]),
    .A2(iX[54]),
    .B1(iX[55]),
    .B2(iY[41]),
    .Y(_02746_));
 sky130_fd_sc_hd__nor2_2 _31178_ (.A(_02745_),
    .B(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__nand2_2 _31179_ (.A(iY[43]),
    .B(iX[53]),
    .Y(_02748_));
 sky130_fd_sc_hd__xnor2_2 _31180_ (.A(_02747_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__o21ba_2 _31181_ (.A1(_02123_),
    .A2(_02125_),
    .B1_N(_02122_),
    .X(_02750_));
 sky130_fd_sc_hd__xnor2_2 _31182_ (.A(_02749_),
    .B(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__and2_2 _31183_ (.A(_02744_),
    .B(_02751_),
    .X(_02753_));
 sky130_fd_sc_hd__nor2_2 _31184_ (.A(_02744_),
    .B(_02751_),
    .Y(_02754_));
 sky130_fd_sc_hd__or2_2 _31185_ (.A(_02753_),
    .B(_02754_),
    .X(_02755_));
 sky130_fd_sc_hd__a21o_2 _31186_ (.A1(_02165_),
    .A2(_02738_),
    .B1(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__nand3_2 _31187_ (.A(_02165_),
    .B(_02738_),
    .C(_02755_),
    .Y(_02757_));
 sky130_fd_sc_hd__o211ai_2 _31188_ (.A1(_02737_),
    .A2(_02130_),
    .B1(_02756_),
    .C1(_02757_),
    .Y(_02758_));
 sky130_fd_sc_hd__a211o_2 _31189_ (.A1(_02756_),
    .A2(_02757_),
    .B1(_02737_),
    .C1(_02130_),
    .X(_02759_));
 sky130_fd_sc_hd__a2bb2o_2 _31190_ (.A1_N(_02735_),
    .A2_N(_02736_),
    .B1(_02758_),
    .B2(_02759_),
    .X(_02760_));
 sky130_fd_sc_hd__and4bb_2 _31191_ (.A_N(_02735_),
    .B_N(_02736_),
    .C(_02758_),
    .D(_02759_),
    .X(_02761_));
 sky130_fd_sc_hd__inv_2 _31192_ (.A(_02761_),
    .Y(_02762_));
 sky130_fd_sc_hd__o211a_2 _31193_ (.A1(_02173_),
    .A2(_02177_),
    .B1(_02760_),
    .C1(_02762_),
    .X(_02764_));
 sky130_fd_sc_hd__a211oi_2 _31194_ (.A1(_02760_),
    .A2(_02762_),
    .B1(_02173_),
    .C1(_02177_),
    .Y(_02765_));
 sky130_fd_sc_hd__inv_2 _31195_ (.A(_02213_),
    .Y(_02766_));
 sky130_fd_sc_hd__and4_2 _31196_ (.A(iX[42]),
    .B(iX[43]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_02767_));
 sky130_fd_sc_hd__a22oi_2 _31197_ (.A1(iX[43]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[42]),
    .Y(_02768_));
 sky130_fd_sc_hd__nor2_2 _31198_ (.A(_02767_),
    .B(_02768_),
    .Y(_02769_));
 sky130_fd_sc_hd__nand2_2 _31199_ (.A(iX[41]),
    .B(iY[55]),
    .Y(_02770_));
 sky130_fd_sc_hd__xnor2_2 _31200_ (.A(_02769_),
    .B(_02770_),
    .Y(_02771_));
 sky130_fd_sc_hd__and4_2 _31201_ (.A(iX[45]),
    .B(iX[46]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_02772_));
 sky130_fd_sc_hd__a22oi_2 _31202_ (.A1(iX[46]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[45]),
    .Y(_02773_));
 sky130_fd_sc_hd__nor2_2 _31203_ (.A(_02772_),
    .B(_02773_),
    .Y(_02775_));
 sky130_fd_sc_hd__nand2_2 _31204_ (.A(iX[44]),
    .B(iY[52]),
    .Y(_02776_));
 sky130_fd_sc_hd__xnor2_2 _31205_ (.A(_02775_),
    .B(_02776_),
    .Y(_02777_));
 sky130_fd_sc_hd__o21ba_2 _31206_ (.A1(_02190_),
    .A2(_02193_),
    .B1_N(_02189_),
    .X(_02778_));
 sky130_fd_sc_hd__xnor2_2 _31207_ (.A(_02777_),
    .B(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__and2_2 _31208_ (.A(_02771_),
    .B(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__nor2_2 _31209_ (.A(_02771_),
    .B(_02779_),
    .Y(_02781_));
 sky130_fd_sc_hd__or2_2 _31210_ (.A(_02780_),
    .B(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__or3_2 _31211_ (.A(_02201_),
    .B(_02206_),
    .C(_02207_),
    .X(_02783_));
 sky130_fd_sc_hd__o21ba_2 _31212_ (.A1(_02118_),
    .A2(_02120_),
    .B1_N(_02117_),
    .X(_02784_));
 sky130_fd_sc_hd__and4_2 _31213_ (.A(iY[47]),
    .B(iX[48]),
    .C(iY[48]),
    .D(iX[49]),
    .X(_02786_));
 sky130_fd_sc_hd__a22oi_2 _31214_ (.A1(iX[48]),
    .A2(iY[48]),
    .B1(iX[49]),
    .B2(iY[47]),
    .Y(_02787_));
 sky130_fd_sc_hd__nand2_2 _31215_ (.A(iX[47]),
    .B(iY[49]),
    .Y(_02788_));
 sky130_fd_sc_hd__o21a_2 _31216_ (.A1(_02786_),
    .A2(_02787_),
    .B1(_02788_),
    .X(_02789_));
 sky130_fd_sc_hd__nor3_2 _31217_ (.A(_02786_),
    .B(_02787_),
    .C(_02788_),
    .Y(_02790_));
 sky130_fd_sc_hd__nor2_2 _31218_ (.A(_02789_),
    .B(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__xnor2_2 _31219_ (.A(_02784_),
    .B(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__o21ai_2 _31220_ (.A1(_02202_),
    .A2(_02207_),
    .B1(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__or3_2 _31221_ (.A(_02202_),
    .B(_02207_),
    .C(_02792_),
    .X(_02794_));
 sky130_fd_sc_hd__nand2_2 _31222_ (.A(_02793_),
    .B(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hd__a21oi_2 _31223_ (.A1(_02783_),
    .A2(_02210_),
    .B1(_02795_),
    .Y(_02797_));
 sky130_fd_sc_hd__and3_2 _31224_ (.A(_02783_),
    .B(_02210_),
    .C(_02795_),
    .X(_02798_));
 sky130_fd_sc_hd__nor3_2 _31225_ (.A(_02782_),
    .B(_02797_),
    .C(_02798_),
    .Y(_02799_));
 sky130_fd_sc_hd__o21a_2 _31226_ (.A1(_02797_),
    .A2(_02798_),
    .B1(_02782_),
    .X(_02800_));
 sky130_fd_sc_hd__a211oi_2 _31227_ (.A1(_02133_),
    .A2(_02135_),
    .B1(_02799_),
    .C1(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__o211a_2 _31228_ (.A1(_02799_),
    .A2(_02800_),
    .B1(_02133_),
    .C1(_02135_),
    .X(_02802_));
 sky130_fd_sc_hd__a211oi_2 _31229_ (.A1(_02766_),
    .A2(_02216_),
    .B1(_02801_),
    .C1(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__o211a_2 _31230_ (.A1(_02801_),
    .A2(_02802_),
    .B1(_02766_),
    .C1(_02216_),
    .X(_02804_));
 sky130_fd_sc_hd__nor4_2 _31231_ (.A(_02764_),
    .B(_02765_),
    .C(_02803_),
    .D(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__o22a_2 _31232_ (.A1(_02764_),
    .A2(_02765_),
    .B1(_02803_),
    .B2(_02804_),
    .X(_02806_));
 sky130_fd_sc_hd__a211o_2 _31233_ (.A1(_02179_),
    .A2(_02223_),
    .B1(_02805_),
    .C1(_02806_),
    .X(_02808_));
 sky130_fd_sc_hd__o211ai_2 _31234_ (.A1(_02805_),
    .A2(_02806_),
    .B1(_02179_),
    .C1(_02223_),
    .Y(_02809_));
 sky130_fd_sc_hd__and2_2 _31235_ (.A(_02808_),
    .B(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__a21bo_2 _31236_ (.A1(_02249_),
    .A2(_02270_),
    .B1_N(_02268_),
    .X(_02811_));
 sky130_fd_sc_hd__or2b_2 _31237_ (.A(_02238_),
    .B_N(_02237_),
    .X(_02812_));
 sky130_fd_sc_hd__and4_2 _31238_ (.A(iX[36]),
    .B(iX[37]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_02813_));
 sky130_fd_sc_hd__a22oi_2 _31239_ (.A1(iX[37]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[36]),
    .Y(_02814_));
 sky130_fd_sc_hd__nor2_2 _31240_ (.A(_02813_),
    .B(_02814_),
    .Y(_02815_));
 sky130_fd_sc_hd__nand2_2 _31241_ (.A(iX[35]),
    .B(iY[61]),
    .Y(_02816_));
 sky130_fd_sc_hd__xnor2_2 _31242_ (.A(_02815_),
    .B(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__o21ba_2 _31243_ (.A1(_02233_),
    .A2(_02235_),
    .B1_N(_02232_),
    .X(_02819_));
 sky130_fd_sc_hd__xnor2_2 _31244_ (.A(_02817_),
    .B(_02819_),
    .Y(_02820_));
 sky130_fd_sc_hd__and2_2 _31245_ (.A(iX[34]),
    .B(iY[62]),
    .X(_02821_));
 sky130_fd_sc_hd__or2_2 _31246_ (.A(_02820_),
    .B(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__nand2_2 _31247_ (.A(_02820_),
    .B(_02821_),
    .Y(_02823_));
 sky130_fd_sc_hd__nand2_2 _31248_ (.A(_02822_),
    .B(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__a21oi_2 _31249_ (.A1(_02812_),
    .A2(_02242_),
    .B1(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__and3_2 _31250_ (.A(_02812_),
    .B(_02242_),
    .C(_02824_),
    .X(_02826_));
 sky130_fd_sc_hd__nor2_2 _31251_ (.A(_02825_),
    .B(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__nand2_2 _31252_ (.A(iX[33]),
    .B(iY[63]),
    .Y(_02828_));
 sky130_fd_sc_hd__xnor2_2 _31253_ (.A(_02827_),
    .B(_02828_),
    .Y(_02830_));
 sky130_fd_sc_hd__or2b_2 _31254_ (.A(_02254_),
    .B_N(_02260_),
    .X(_02831_));
 sky130_fd_sc_hd__or2b_2 _31255_ (.A(_02253_),
    .B_N(_02261_),
    .X(_02832_));
 sky130_fd_sc_hd__and2b_2 _31256_ (.A_N(_02195_),
    .B(_02194_),
    .X(_02833_));
 sky130_fd_sc_hd__o21ba_2 _31257_ (.A1(_02256_),
    .A2(_02259_),
    .B1_N(_02255_),
    .X(_02834_));
 sky130_fd_sc_hd__o21ba_2 _31258_ (.A1(_02185_),
    .A2(_02187_),
    .B1_N(_02184_),
    .X(_02835_));
 sky130_fd_sc_hd__and4_2 _31259_ (.A(iX[39]),
    .B(iX[40]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_02836_));
 sky130_fd_sc_hd__a22oi_2 _31260_ (.A1(iX[40]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[39]),
    .Y(_02837_));
 sky130_fd_sc_hd__nor2_2 _31261_ (.A(_02836_),
    .B(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__nand2_2 _31262_ (.A(iX[38]),
    .B(iY[58]),
    .Y(_02839_));
 sky130_fd_sc_hd__xnor2_2 _31263_ (.A(_02838_),
    .B(_02839_),
    .Y(_02841_));
 sky130_fd_sc_hd__xnor2_2 _31264_ (.A(_02835_),
    .B(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__xnor2_2 _31265_ (.A(_02834_),
    .B(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__o21a_2 _31266_ (.A1(_02833_),
    .A2(_02197_),
    .B1(_02843_),
    .X(_02844_));
 sky130_fd_sc_hd__nor3_2 _31267_ (.A(_02833_),
    .B(_02197_),
    .C(_02843_),
    .Y(_02845_));
 sky130_fd_sc_hd__a211oi_2 _31268_ (.A1(_02831_),
    .A2(_02832_),
    .B1(_02844_),
    .C1(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__o211a_2 _31269_ (.A1(_02844_),
    .A2(_02845_),
    .B1(_02831_),
    .C1(_02832_),
    .X(_02847_));
 sky130_fd_sc_hd__nor2_2 _31270_ (.A(_02263_),
    .B(_02265_),
    .Y(_02848_));
 sky130_fd_sc_hd__or3_2 _31271_ (.A(_02846_),
    .B(_02847_),
    .C(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__o21ai_2 _31272_ (.A1(_02846_),
    .A2(_02847_),
    .B1(_02848_),
    .Y(_02850_));
 sky130_fd_sc_hd__and3_2 _31273_ (.A(_02830_),
    .B(_02849_),
    .C(_02850_),
    .X(_02852_));
 sky130_fd_sc_hd__a21oi_2 _31274_ (.A1(_02849_),
    .A2(_02850_),
    .B1(_02830_),
    .Y(_02853_));
 sky130_fd_sc_hd__nor2_2 _31275_ (.A(_02852_),
    .B(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hd__o21a_2 _31276_ (.A1(_02219_),
    .A2(_02221_),
    .B1(_02854_),
    .X(_02855_));
 sky130_fd_sc_hd__nor2_2 _31277_ (.A(_02219_),
    .B(_02221_),
    .Y(_02856_));
 sky130_fd_sc_hd__and2b_2 _31278_ (.A_N(_02854_),
    .B(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__or2_2 _31279_ (.A(_02855_),
    .B(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__xnor2_2 _31280_ (.A(_02811_),
    .B(_02858_),
    .Y(_02859_));
 sky130_fd_sc_hd__nand2_2 _31281_ (.A(_02810_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__or2_2 _31282_ (.A(_02810_),
    .B(_02859_),
    .X(_02861_));
 sky130_fd_sc_hd__nand2_2 _31283_ (.A(_02860_),
    .B(_02861_),
    .Y(_02863_));
 sky130_fd_sc_hd__inv_2 _31284_ (.A(_02227_),
    .Y(_02864_));
 sky130_fd_sc_hd__o31a_2 _31285_ (.A1(_02229_),
    .A2(_02276_),
    .A3(_02277_),
    .B1(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__or2_2 _31286_ (.A(_02863_),
    .B(_02865_),
    .X(_02866_));
 sky130_fd_sc_hd__nand2_2 _31287_ (.A(_02863_),
    .B(_02865_),
    .Y(_02867_));
 sky130_fd_sc_hd__nand2_2 _31288_ (.A(_02866_),
    .B(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__nor2_2 _31289_ (.A(_02274_),
    .B(_02276_),
    .Y(_02869_));
 sky130_fd_sc_hd__or2_2 _31290_ (.A(_02868_),
    .B(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__nand2_2 _31291_ (.A(_02868_),
    .B(_02869_),
    .Y(_02871_));
 sky130_fd_sc_hd__nand2_2 _31292_ (.A(_02870_),
    .B(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__and2_2 _31293_ (.A(_02281_),
    .B(_02283_),
    .X(_02874_));
 sky130_fd_sc_hd__or2_2 _31294_ (.A(_02872_),
    .B(_02874_),
    .X(_02875_));
 sky130_fd_sc_hd__nand2_2 _31295_ (.A(_02872_),
    .B(_02874_),
    .Y(_02876_));
 sky130_fd_sc_hd__and2_2 _31296_ (.A(_02875_),
    .B(_02876_),
    .X(_02877_));
 sky130_fd_sc_hd__nand2b_2 _31297_ (.A_N(_02701_),
    .B(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__or2b_2 _31298_ (.A(_02877_),
    .B_N(_02701_),
    .X(_02879_));
 sky130_fd_sc_hd__a21oi_2 _31299_ (.A1(_02046_),
    .A2(_02289_),
    .B1(_02287_),
    .Y(_02880_));
 sky130_fd_sc_hd__inv_2 _31300_ (.A(_02880_),
    .Y(_02881_));
 sky130_fd_sc_hd__and3_2 _31301_ (.A(_02878_),
    .B(_02879_),
    .C(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__a21oi_2 _31302_ (.A1(_02878_),
    .A2(_02879_),
    .B1(_02881_),
    .Y(_02883_));
 sky130_fd_sc_hd__or2_2 _31303_ (.A(_02882_),
    .B(_02883_),
    .X(_02885_));
 sky130_fd_sc_hd__a21oi_2 _31304_ (.A1(_02699_),
    .A2(_02700_),
    .B1(_02885_),
    .Y(_02886_));
 sky130_fd_sc_hd__and3_2 _31305_ (.A(_02699_),
    .B(_02700_),
    .C(_02885_),
    .X(_02887_));
 sky130_fd_sc_hd__nor2_2 _31306_ (.A(_02886_),
    .B(_02887_),
    .Y(_02888_));
 sky130_fd_sc_hd__xor2_2 _31307_ (.A(_02698_),
    .B(_02888_),
    .X(_02889_));
 sky130_fd_sc_hd__nand2_2 _31308_ (.A(_11370_),
    .B(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__or2_2 _31309_ (.A(_11370_),
    .B(_02889_),
    .X(_02891_));
 sky130_fd_sc_hd__nand2_2 _31310_ (.A(_02890_),
    .B(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__inv_2 _31311_ (.A(oO[31]),
    .Y(_02893_));
 sky130_fd_sc_hd__inv_2 _31312_ (.A(_02294_),
    .Y(_02894_));
 sky130_fd_sc_hd__nor2_2 _31313_ (.A(_02894_),
    .B(_02498_),
    .Y(_02896_));
 sky130_fd_sc_hd__a21oi_2 _31314_ (.A1(_02893_),
    .A2(_02499_),
    .B1(_02896_),
    .Y(_02897_));
 sky130_fd_sc_hd__or2_2 _31315_ (.A(_02892_),
    .B(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__nand2_2 _31316_ (.A(_02892_),
    .B(_02897_),
    .Y(_02899_));
 sky130_fd_sc_hd__nand2_2 _31317_ (.A(_02898_),
    .B(_02899_),
    .Y(_02900_));
 sky130_fd_sc_hd__nand2_2 _31318_ (.A(_02113_),
    .B(_02501_),
    .Y(_02901_));
 sky130_fd_sc_hd__a21o_2 _31319_ (.A1(_02111_),
    .A2(_02101_),
    .B1(_02502_),
    .X(_02902_));
 sky130_fd_sc_hd__and2_2 _31320_ (.A(_02901_),
    .B(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__xnor2_2 _31321_ (.A(_02900_),
    .B(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__or2_2 _31322_ (.A(_11383_),
    .B(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__nand2_2 _31323_ (.A(_11383_),
    .B(_02904_),
    .Y(_02907_));
 sky130_fd_sc_hd__nand2_2 _31324_ (.A(_02905_),
    .B(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__a21boi_2 _31325_ (.A1(_02510_),
    .A2(_02107_),
    .B1_N(_02509_),
    .Y(_02909_));
 sky130_fd_sc_hd__nor2_2 _31326_ (.A(_02507_),
    .B(_02909_),
    .Y(_02910_));
 sky130_fd_sc_hd__xor2_2 _31327_ (.A(_02908_),
    .B(_02910_),
    .X(oO[64]));
 sky130_fd_sc_hd__or2_2 _31328_ (.A(_02698_),
    .B(_02888_),
    .X(_02911_));
 sky130_fd_sc_hd__nand2_2 _31329_ (.A(_11560_),
    .B(_11561_),
    .Y(_02912_));
 sky130_fd_sc_hd__or2b_2 _31330_ (.A(_02688_),
    .B_N(_02687_),
    .X(_02913_));
 sky130_fd_sc_hd__nand2_2 _31331_ (.A(_02513_),
    .B(_02689_),
    .Y(_02914_));
 sky130_fd_sc_hd__and2_2 _31332_ (.A(_02519_),
    .B(_02556_),
    .X(_02915_));
 sky130_fd_sc_hd__and2b_2 _31333_ (.A_N(_02557_),
    .B(_02517_),
    .X(_02917_));
 sky130_fd_sc_hd__inv_2 _31334_ (.A(_02325_),
    .Y(_02918_));
 sky130_fd_sc_hd__o2bb2a_2 _31335_ (.A1_N(_02918_),
    .A2_N(_02537_),
    .B1(_02536_),
    .B2(_02535_),
    .X(_02919_));
 sky130_fd_sc_hd__o21ba_2 _31336_ (.A1(_02915_),
    .A2(_02917_),
    .B1_N(_02919_),
    .X(_02920_));
 sky130_fd_sc_hd__or3b_2 _31337_ (.A(_02915_),
    .B(_02917_),
    .C_N(_02919_),
    .X(_02921_));
 sky130_fd_sc_hd__and2b_2 _31338_ (.A_N(_02920_),
    .B(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__nand2_2 _31339_ (.A(_02552_),
    .B(_02553_),
    .Y(_02923_));
 sky130_fd_sc_hd__nor2_2 _31340_ (.A(_02552_),
    .B(_02553_),
    .Y(_02924_));
 sky130_fd_sc_hd__a21o_2 _31341_ (.A1(_02538_),
    .A2(_02923_),
    .B1(_02924_),
    .X(_02925_));
 sky130_fd_sc_hd__or2b_2 _31342_ (.A(_02599_),
    .B_N(_02601_),
    .X(_02926_));
 sky130_fd_sc_hd__buf_1 _31343_ (.A(_01522_),
    .X(_02928_));
 sky130_fd_sc_hd__and2_2 _31344_ (.A(_02529_),
    .B(_02533_),
    .X(_02929_));
 sky130_fd_sc_hd__a31o_2 _31345_ (.A1(_18749_),
    .A2(_02928_),
    .A3(_02531_),
    .B1(_02929_),
    .X(_02930_));
 sky130_fd_sc_hd__or4b_2 _31346_ (.A(_18120_),
    .B(_16271_),
    .C(_01746_),
    .D_N(_01521_),
    .X(_02931_));
 sky130_fd_sc_hd__a2bb2o_2 _31347_ (.A1_N(_18120_),
    .A2_N(_01746_),
    .B1(_01521_),
    .B2(_14629_),
    .X(_02932_));
 sky130_fd_sc_hd__nand2_2 _31348_ (.A(_02931_),
    .B(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__nor2_2 _31349_ (.A(_16625_),
    .B(_02322_),
    .Y(_02934_));
 sky130_fd_sc_hd__xor2_2 _31350_ (.A(_02933_),
    .B(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__and4_2 _31351_ (.A(_16268_),
    .B(_16277_),
    .C(_00161_),
    .D(_00564_),
    .X(_02936_));
 sky130_fd_sc_hd__a22o_2 _31352_ (.A1(_02338_),
    .A2(_00161_),
    .B1(_00565_),
    .B2(_01564_),
    .X(_02937_));
 sky130_fd_sc_hd__or4b_2 _31353_ (.A(_18368_),
    .B(_00943_),
    .C(_02936_),
    .D_N(_02937_),
    .X(_02939_));
 sky130_fd_sc_hd__xor2_2 _31354_ (.A(_00157_),
    .B(_00160_),
    .X(_02940_));
 sky130_fd_sc_hd__or4_2 _31355_ (.A(_00195_),
    .B(_00589_),
    .C(_02940_),
    .D(_01512_),
    .X(_02941_));
 sky130_fd_sc_hd__a22o_2 _31356_ (.A1(_18754_),
    .A2(_01510_),
    .B1(_02941_),
    .B2(_02937_),
    .X(_02942_));
 sky130_fd_sc_hd__a31o_2 _31357_ (.A1(_14629_),
    .A2(_01510_),
    .A3(_02523_),
    .B1(_02522_),
    .X(_02943_));
 sky130_fd_sc_hd__and3_2 _31358_ (.A(_02939_),
    .B(_02942_),
    .C(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__a21oi_2 _31359_ (.A1(_02939_),
    .A2(_02942_),
    .B1(_02943_),
    .Y(_02945_));
 sky130_fd_sc_hd__nor2_2 _31360_ (.A(_02944_),
    .B(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__xor2_2 _31361_ (.A(_02935_),
    .B(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__and2b_2 _31362_ (.A_N(_02527_),
    .B(_02525_),
    .X(_02948_));
 sky130_fd_sc_hd__a21o_2 _31363_ (.A1(_02528_),
    .A2(_02534_),
    .B1(_02948_),
    .X(_02950_));
 sky130_fd_sc_hd__xnor2_2 _31364_ (.A(_02947_),
    .B(_02950_),
    .Y(_02951_));
 sky130_fd_sc_hd__xnor2_2 _31365_ (.A(_02930_),
    .B(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__or2b_2 _31366_ (.A(_02542_),
    .B_N(_02548_),
    .X(_02953_));
 sky130_fd_sc_hd__a21bo_2 _31367_ (.A1(_02541_),
    .A2(_02549_),
    .B1_N(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__a21o_2 _31368_ (.A1(_02568_),
    .A2(_02578_),
    .B1(_02577_),
    .X(_02955_));
 sky130_fd_sc_hd__buf_1 _31369_ (.A(_18729_),
    .X(_02956_));
 sky130_fd_sc_hd__nor2_2 _31370_ (.A(_02545_),
    .B(_02546_),
    .Y(_02957_));
 sky130_fd_sc_hd__a31o_2 _31371_ (.A1(_02338_),
    .A2(_02956_),
    .A3(_02547_),
    .B1(_02957_),
    .X(_02958_));
 sky130_fd_sc_hd__a21bo_2 _31372_ (.A1(_02562_),
    .A2(_02566_),
    .B1_N(_02564_),
    .X(_02959_));
 sky130_fd_sc_hd__nand2_2 _31373_ (.A(_14648_),
    .B(_18732_),
    .Y(_02961_));
 sky130_fd_sc_hd__or3_4 _31374_ (.A(_15211_),
    .B(_18110_),
    .C(_18112_),
    .X(_02962_));
 sky130_fd_sc_hd__xor2_2 _31375_ (.A(_02961_),
    .B(_02962_),
    .X(_02963_));
 sky130_fd_sc_hd__nand2_2 _31376_ (.A(_01784_),
    .B(_18729_),
    .Y(_02964_));
 sky130_fd_sc_hd__xor2_2 _31377_ (.A(_02963_),
    .B(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__xnor2_2 _31378_ (.A(_02959_),
    .B(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__xnor2_2 _31379_ (.A(_02958_),
    .B(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__xnor2_2 _31380_ (.A(_02955_),
    .B(_02967_),
    .Y(_02968_));
 sky130_fd_sc_hd__xnor2_2 _31381_ (.A(_02954_),
    .B(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__and2_2 _31382_ (.A(_02540_),
    .B(_02550_),
    .X(_02970_));
 sky130_fd_sc_hd__a21oi_2 _31383_ (.A1(_02539_),
    .A2(_02551_),
    .B1(_02970_),
    .Y(_02972_));
 sky130_fd_sc_hd__xor2_2 _31384_ (.A(_02969_),
    .B(_02972_),
    .X(_02973_));
 sky130_fd_sc_hd__xnor2_2 _31385_ (.A(_02952_),
    .B(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__xnor2_2 _31386_ (.A(_02926_),
    .B(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__xor2_2 _31387_ (.A(_02925_),
    .B(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__or2_2 _31388_ (.A(_02592_),
    .B(_02595_),
    .X(_02977_));
 sky130_fd_sc_hd__o21ai_2 _31389_ (.A1(_02580_),
    .A2(_02596_),
    .B1(_02977_),
    .Y(_02978_));
 sky130_fd_sc_hd__or2b_2 _31390_ (.A(_02623_),
    .B_N(_02606_),
    .X(_02979_));
 sky130_fd_sc_hd__or2b_2 _31391_ (.A(_02605_),
    .B_N(_02624_),
    .X(_02980_));
 sky130_fd_sc_hd__or3_2 _31392_ (.A(_15005_),
    .B(_17408_),
    .C(_02563_),
    .X(_02981_));
 sky130_fd_sc_hd__buf_1 _31393_ (.A(_16292_),
    .X(_02983_));
 sky130_fd_sc_hd__buf_1 _31394_ (.A(_17630_),
    .X(_02984_));
 sky130_fd_sc_hd__a22o_2 _31395_ (.A1(_02983_),
    .A2(_17394_),
    .B1(_02984_),
    .B2(_15888_),
    .X(_02985_));
 sky130_fd_sc_hd__and2_2 _31396_ (.A(_02981_),
    .B(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__nor2_2 _31397_ (.A(_01576_),
    .B(_17628_),
    .Y(_02987_));
 sky130_fd_sc_hd__xnor2_2 _31398_ (.A(_02986_),
    .B(_02987_),
    .Y(_02988_));
 sky130_fd_sc_hd__buf_1 _31399_ (.A(_17460_),
    .X(_02989_));
 sky130_fd_sc_hd__nor2_2 _31400_ (.A(_16312_),
    .B(_16258_),
    .Y(_02990_));
 sky130_fd_sc_hd__o22a_2 _31401_ (.A1(_01832_),
    .A2(_00996_),
    .B1(_16258_),
    .B2(_18181_),
    .X(_02991_));
 sky130_fd_sc_hd__a31o_2 _31402_ (.A1(_02989_),
    .A2(_16934_),
    .A3(_02990_),
    .B1(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__buf_1 _31403_ (.A(_15679_),
    .X(_02994_));
 sky130_fd_sc_hd__nand2_2 _31404_ (.A(_02994_),
    .B(_16614_),
    .Y(_02995_));
 sky130_fd_sc_hd__xnor2_2 _31405_ (.A(_02992_),
    .B(_02995_),
    .Y(_02996_));
 sky130_fd_sc_hd__a21o_2 _31406_ (.A1(_02569_),
    .A2(_02573_),
    .B1(_02571_),
    .X(_02997_));
 sky130_fd_sc_hd__xor2_2 _31407_ (.A(_02996_),
    .B(_02997_),
    .X(_02998_));
 sky130_fd_sc_hd__xor2_2 _31408_ (.A(_02988_),
    .B(_02998_),
    .X(_02999_));
 sky130_fd_sc_hd__or2b_2 _31409_ (.A(_02468_),
    .B_N(_02586_),
    .X(_03000_));
 sky130_fd_sc_hd__a31o_2 _31410_ (.A1(_14606_),
    .A2(_01837_),
    .A3(_02611_),
    .B1(_02607_),
    .X(_03001_));
 sky130_fd_sc_hd__nor2_2 _31411_ (.A(_15154_),
    .B(_00255_),
    .Y(_03002_));
 sky130_fd_sc_hd__nor2_2 _31412_ (.A(_14948_),
    .B(_17007_),
    .Y(_03003_));
 sky130_fd_sc_hd__xnor2_2 _31413_ (.A(_03002_),
    .B(_03003_),
    .Y(_03005_));
 sky130_fd_sc_hd__nor2_2 _31414_ (.A(_15598_),
    .B(_01828_),
    .Y(_03006_));
 sky130_fd_sc_hd__xnor2_2 _31415_ (.A(_03005_),
    .B(_03006_),
    .Y(_03007_));
 sky130_fd_sc_hd__xnor2_2 _31416_ (.A(_03001_),
    .B(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__a21oi_2 _31417_ (.A1(_02584_),
    .A2(_03000_),
    .B1(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__and3_2 _31418_ (.A(_02584_),
    .B(_03000_),
    .C(_03008_),
    .X(_03010_));
 sky130_fd_sc_hd__or2_2 _31419_ (.A(_03009_),
    .B(_03010_),
    .X(_03011_));
 sky130_fd_sc_hd__a21oi_2 _31420_ (.A1(_02581_),
    .A2(_02591_),
    .B1(_02589_),
    .Y(_03012_));
 sky130_fd_sc_hd__xor2_2 _31421_ (.A(_03011_),
    .B(_03012_),
    .X(_03013_));
 sky130_fd_sc_hd__and2_2 _31422_ (.A(_02999_),
    .B(_03013_),
    .X(_03014_));
 sky130_fd_sc_hd__nor2_2 _31423_ (.A(_02999_),
    .B(_03013_),
    .Y(_03016_));
 sky130_fd_sc_hd__a211oi_2 _31424_ (.A1(_02979_),
    .A2(_02980_),
    .B1(_03014_),
    .C1(_03016_),
    .Y(_03017_));
 sky130_fd_sc_hd__o211a_2 _31425_ (.A1(_03014_),
    .A2(_03016_),
    .B1(_02979_),
    .C1(_02980_),
    .X(_03018_));
 sky130_fd_sc_hd__nor2_2 _31426_ (.A(_03017_),
    .B(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hd__xor2_2 _31427_ (.A(_02978_),
    .B(_03019_),
    .X(_03020_));
 sky130_fd_sc_hd__a32oi_2 _31428_ (.A1(_02617_),
    .A2(_02618_),
    .A3(_02621_),
    .B1(_02622_),
    .B2(_02612_),
    .Y(_03021_));
 sky130_fd_sc_hd__a21oi_2 _31429_ (.A1(_02628_),
    .A2(_02638_),
    .B1(_02637_),
    .Y(_03022_));
 sky130_fd_sc_hd__buf_1 _31430_ (.A(_14606_),
    .X(_03023_));
 sky130_fd_sc_hd__buf_1 _31431_ (.A(_17702_),
    .X(_03024_));
 sky130_fd_sc_hd__and4_2 _31432_ (.A(_01039_),
    .B(_14411_),
    .C(_18209_),
    .D(_18463_),
    .X(_03025_));
 sky130_fd_sc_hd__o22a_2 _31433_ (.A1(_01605_),
    .A2(_18200_),
    .B1(_18443_),
    .B2(_02608_),
    .X(_03027_));
 sky130_fd_sc_hd__nor2_2 _31434_ (.A(_03025_),
    .B(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__a21oi_2 _31435_ (.A1(_03023_),
    .A2(_03024_),
    .B1(_03028_),
    .Y(_03029_));
 sky130_fd_sc_hd__and3_2 _31436_ (.A(_14606_),
    .B(_03024_),
    .C(_03028_),
    .X(_03030_));
 sky130_fd_sc_hd__nor2_2 _31437_ (.A(_03029_),
    .B(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__or4_2 _31438_ (.A(_14625_),
    .B(_18791_),
    .C(_00271_),
    .D(_00666_),
    .X(_03032_));
 sky130_fd_sc_hd__a22o_2 _31439_ (.A1(_13544_),
    .A2(_01647_),
    .B1(_00268_),
    .B2(_17463_),
    .X(_03033_));
 sky130_fd_sc_hd__nand2_2 _31440_ (.A(_03032_),
    .B(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__nand2_2 _31441_ (.A(_13889_),
    .B(_00662_),
    .Y(_03035_));
 sky130_fd_sc_hd__xnor2_2 _31442_ (.A(_03034_),
    .B(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__a21oi_2 _31443_ (.A1(_02614_),
    .A2(_02617_),
    .B1(_03036_),
    .Y(_03038_));
 sky130_fd_sc_hd__and3_2 _31444_ (.A(_02614_),
    .B(_02617_),
    .C(_03036_),
    .X(_03039_));
 sky130_fd_sc_hd__or2_2 _31445_ (.A(_03038_),
    .B(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__xnor2_2 _31446_ (.A(_03031_),
    .B(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__xnor2_2 _31447_ (.A(_03022_),
    .B(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__xnor2_2 _31448_ (.A(_03021_),
    .B(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__a31o_2 _31449_ (.A1(_02626_),
    .A2(_01862_),
    .A3(_02634_),
    .B1(_02633_),
    .X(_03044_));
 sky130_fd_sc_hd__nand2_2 _31450_ (.A(_02626_),
    .B(_02629_),
    .Y(_03045_));
 sky130_fd_sc_hd__nor2_2 _31451_ (.A(_12848_),
    .B(_01087_),
    .Y(_03046_));
 sky130_fd_sc_hd__and3_2 _31452_ (.A(_15887_),
    .B(_01650_),
    .C(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__o22a_2 _31453_ (.A1(_12848_),
    .A2(_01866_),
    .B1(_02647_),
    .B2(_15646_),
    .X(_03049_));
 sky130_fd_sc_hd__nor2_2 _31454_ (.A(_03047_),
    .B(_03049_),
    .Y(_03050_));
 sky130_fd_sc_hd__xnor2_2 _31455_ (.A(_03045_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__o21ai_2 _31456_ (.A1(_02645_),
    .A2(_02649_),
    .B1(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__or3_2 _31457_ (.A(_02645_),
    .B(_02649_),
    .C(_03051_),
    .X(_03053_));
 sky130_fd_sc_hd__and3_2 _31458_ (.A(_03044_),
    .B(_03052_),
    .C(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__a21oi_2 _31459_ (.A1(_03052_),
    .A2(_03053_),
    .B1(_03044_),
    .Y(_03055_));
 sky130_fd_sc_hd__nor2_2 _31460_ (.A(_03054_),
    .B(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__nor2_2 _31461_ (.A(_14978_),
    .B(_02391_),
    .Y(_03057_));
 sky130_fd_sc_hd__or3_2 _31462_ (.A(_11794_),
    .B(_02397_),
    .C(_02398_),
    .X(_03058_));
 sky130_fd_sc_hd__xnor2_2 _31463_ (.A(_02644_),
    .B(_03058_),
    .Y(_03060_));
 sky130_fd_sc_hd__xor2_2 _31464_ (.A(_03057_),
    .B(_03060_),
    .X(_03061_));
 sky130_fd_sc_hd__inv_2 _31465_ (.A(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__and2_2 _31466_ (.A(_02658_),
    .B(_02660_),
    .X(_03063_));
 sky130_fd_sc_hd__nor2_2 _31467_ (.A(_03063_),
    .B(_02663_),
    .Y(_03064_));
 sky130_fd_sc_hd__o22a_2 _31468_ (.A1(_11571_),
    .A2(_03063_),
    .B1(_02663_),
    .B2(_11576_),
    .X(_03065_));
 sky130_fd_sc_hd__a31o_2 _31469_ (.A1(_17392_),
    .A2(_11585_),
    .A3(_03064_),
    .B1(_03065_),
    .X(_03066_));
 sky130_fd_sc_hd__a21o_2 _31470_ (.A1(_02658_),
    .A2(_02660_),
    .B1(_02663_),
    .X(_03067_));
 sky130_fd_sc_hd__buf_1 _31471_ (.A(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__a2bb2oi_2 _31472_ (.A1_N(_11382_),
    .A2_N(_03068_),
    .B1(_02666_),
    .B2(_02654_),
    .Y(_03069_));
 sky130_fd_sc_hd__xnor2_2 _31473_ (.A(_03066_),
    .B(_03069_),
    .Y(_03071_));
 sky130_fd_sc_hd__xnor2_2 _31474_ (.A(_03062_),
    .B(_03071_),
    .Y(_03072_));
 sky130_fd_sc_hd__and2b_2 _31475_ (.A_N(_02667_),
    .B(_02668_),
    .X(_03073_));
 sky130_fd_sc_hd__or2b_2 _31476_ (.A(_02668_),
    .B_N(_02667_),
    .X(_03074_));
 sky130_fd_sc_hd__o21a_2 _31477_ (.A1(_02651_),
    .A2(_03073_),
    .B1(_03074_),
    .X(_03075_));
 sky130_fd_sc_hd__xor2_2 _31478_ (.A(_03072_),
    .B(_03075_),
    .X(_03076_));
 sky130_fd_sc_hd__xor2_2 _31479_ (.A(_03056_),
    .B(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__nor2_2 _31480_ (.A(_02670_),
    .B(_02671_),
    .Y(_03078_));
 sky130_fd_sc_hd__nand2_2 _31481_ (.A(_02670_),
    .B(_02671_),
    .Y(_03079_));
 sky130_fd_sc_hd__o21a_2 _31482_ (.A1(_02640_),
    .A2(_03078_),
    .B1(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__xnor2_2 _31483_ (.A(_03077_),
    .B(_03080_),
    .Y(_03082_));
 sky130_fd_sc_hd__xnor2_2 _31484_ (.A(_03043_),
    .B(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__and2b_2 _31485_ (.A_N(_02674_),
    .B(_02673_),
    .X(_03084_));
 sky130_fd_sc_hd__a21oi_2 _31486_ (.A1(_02625_),
    .A2(_02676_),
    .B1(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__xor2_2 _31487_ (.A(_03083_),
    .B(_03085_),
    .X(_03086_));
 sky130_fd_sc_hd__xor2_2 _31488_ (.A(_03020_),
    .B(_03086_),
    .X(_03087_));
 sky130_fd_sc_hd__and2b_2 _31489_ (.A_N(_02677_),
    .B(_02678_),
    .X(_03088_));
 sky130_fd_sc_hd__a21oi_2 _31490_ (.A1(_02603_),
    .A2(_02679_),
    .B1(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__xor2_2 _31491_ (.A(_03087_),
    .B(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__xnor2_2 _31492_ (.A(_02976_),
    .B(_03090_),
    .Y(_03091_));
 sky130_fd_sc_hd__and2b_2 _31493_ (.A_N(_02681_),
    .B(_02680_),
    .X(_03093_));
 sky130_fd_sc_hd__a21oi_2 _31494_ (.A1(_02558_),
    .A2(_02682_),
    .B1(_03093_),
    .Y(_03094_));
 sky130_fd_sc_hd__xor2_2 _31495_ (.A(_03091_),
    .B(_03094_),
    .X(_03095_));
 sky130_fd_sc_hd__xnor2_2 _31496_ (.A(_02922_),
    .B(_03095_),
    .Y(_03096_));
 sky130_fd_sc_hd__and2b_2 _31497_ (.A_N(_02683_),
    .B(_02684_),
    .X(_03097_));
 sky130_fd_sc_hd__a21oi_2 _31498_ (.A1(_02516_),
    .A2(_02685_),
    .B1(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__xor2_2 _31499_ (.A(_03096_),
    .B(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__xnor2_2 _31500_ (.A(_02514_),
    .B(_03099_),
    .Y(_03100_));
 sky130_fd_sc_hd__a21oi_2 _31501_ (.A1(_02913_),
    .A2(_02914_),
    .B1(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__and3_2 _31502_ (.A(_02913_),
    .B(_02914_),
    .C(_03100_),
    .X(_03102_));
 sky130_fd_sc_hd__or2_2 _31503_ (.A(_03101_),
    .B(_03102_),
    .X(_03104_));
 sky130_fd_sc_hd__nand3_2 _31504_ (.A(_01126_),
    .B(_01131_),
    .C(_02693_),
    .Y(_03105_));
 sky130_fd_sc_hd__nand2_2 _31505_ (.A(_02693_),
    .B(_02694_),
    .Y(_03106_));
 sky130_fd_sc_hd__or2b_2 _31506_ (.A(_02493_),
    .B_N(_02690_),
    .X(_03107_));
 sky130_fd_sc_hd__inv_2 _31507_ (.A(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__a31o_2 _31508_ (.A1(_02691_),
    .A2(_03105_),
    .A3(_03106_),
    .B1(_03108_),
    .X(_03109_));
 sky130_fd_sc_hd__xnor2_2 _31509_ (.A(_03104_),
    .B(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__a22oi_2 _31510_ (.A1(iY[35]),
    .A2(iX[62]),
    .B1(iX[63]),
    .B2(iY[34]),
    .Y(_03111_));
 sky130_fd_sc_hd__a31oi_2 _31511_ (.A1(iY[35]),
    .A2(iX[63]),
    .A3(_02704_),
    .B1(_03111_),
    .Y(_03112_));
 sky130_fd_sc_hd__a31o_2 _31512_ (.A1(iY[33]),
    .A2(iX[63]),
    .A3(_02706_),
    .B1(_02705_),
    .X(_03113_));
 sky130_fd_sc_hd__xor2_2 _31513_ (.A(_03112_),
    .B(_03113_),
    .X(_03115_));
 sky130_fd_sc_hd__a21oi_2 _31514_ (.A1(iY[37]),
    .A2(iX[60]),
    .B1(_01373_),
    .Y(_03116_));
 sky130_fd_sc_hd__and3_2 _31515_ (.A(iY[37]),
    .B(iX[60]),
    .C(_01373_),
    .X(_03117_));
 sky130_fd_sc_hd__nor2_2 _31516_ (.A(_03116_),
    .B(_03117_),
    .Y(_03118_));
 sky130_fd_sc_hd__xnor2_2 _31517_ (.A(_03115_),
    .B(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__or2b_2 _31518_ (.A(_02711_),
    .B_N(_02710_),
    .X(_03120_));
 sky130_fd_sc_hd__o21a_2 _31519_ (.A1(_02712_),
    .A2(_02715_),
    .B1(_03120_),
    .X(_03121_));
 sky130_fd_sc_hd__xnor2_2 _31520_ (.A(_03119_),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__a31o_2 _31521_ (.A1(iY[40]),
    .A2(iX[56]),
    .A3(_02725_),
    .B1(_02724_),
    .X(_03123_));
 sky130_fd_sc_hd__nand2_2 _31522_ (.A(iY[38]),
    .B(iX[59]),
    .Y(_03124_));
 sky130_fd_sc_hd__nand2_2 _31523_ (.A(iY[39]),
    .B(iX[59]),
    .Y(_03125_));
 sky130_fd_sc_hd__nor2_2 _31524_ (.A(_02722_),
    .B(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__a21oi_2 _31525_ (.A1(_02723_),
    .A2(_03124_),
    .B1(_03126_),
    .Y(_03127_));
 sky130_fd_sc_hd__nand2_2 _31526_ (.A(iY[40]),
    .B(iX[57]),
    .Y(_03128_));
 sky130_fd_sc_hd__xnor2_2 _31527_ (.A(_03127_),
    .B(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__nand2_2 _31528_ (.A(_02714_),
    .B(_03129_),
    .Y(_03130_));
 sky130_fd_sc_hd__or2_2 _31529_ (.A(_02714_),
    .B(_03129_),
    .X(_03131_));
 sky130_fd_sc_hd__nand2_2 _31530_ (.A(_03130_),
    .B(_03131_),
    .Y(_03132_));
 sky130_fd_sc_hd__xor2_2 _31531_ (.A(_03123_),
    .B(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__nor2_2 _31532_ (.A(_03122_),
    .B(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__and2_2 _31533_ (.A(_03122_),
    .B(_03133_),
    .X(_03136_));
 sky130_fd_sc_hd__nor2_2 _31534_ (.A(_03134_),
    .B(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__o21ai_2 _31535_ (.A1(_02717_),
    .A2(_02733_),
    .B1(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__or3_2 _31536_ (.A(_02717_),
    .B(_02733_),
    .C(_03137_),
    .X(_03139_));
 sky130_fd_sc_hd__and2_2 _31537_ (.A(_03138_),
    .B(_03139_),
    .X(_03140_));
 sky130_fd_sc_hd__and2b_2 _31538_ (.A_N(_02750_),
    .B(_02749_),
    .X(_03141_));
 sky130_fd_sc_hd__nand2_2 _31539_ (.A(_02720_),
    .B(_02731_),
    .Y(_03142_));
 sky130_fd_sc_hd__and4_2 _31540_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[52]),
    .D(iX[53]),
    .X(_03143_));
 sky130_fd_sc_hd__a22oi_2 _31541_ (.A1(iY[45]),
    .A2(iX[52]),
    .B1(iX[53]),
    .B2(iY[44]),
    .Y(_03144_));
 sky130_fd_sc_hd__nor2_2 _31542_ (.A(_03143_),
    .B(_03144_),
    .Y(_03145_));
 sky130_fd_sc_hd__nand2_2 _31543_ (.A(iY[46]),
    .B(iX[51]),
    .Y(_03147_));
 sky130_fd_sc_hd__xnor2_2 _31544_ (.A(_03145_),
    .B(_03147_),
    .Y(_03148_));
 sky130_fd_sc_hd__and4_2 _31545_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[55]),
    .D(iX[56]),
    .X(_03149_));
 sky130_fd_sc_hd__a22oi_2 _31546_ (.A1(iY[42]),
    .A2(iX[55]),
    .B1(iX[56]),
    .B2(iY[41]),
    .Y(_03150_));
 sky130_fd_sc_hd__nor2_2 _31547_ (.A(_03149_),
    .B(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__nand2_2 _31548_ (.A(iY[43]),
    .B(iX[54]),
    .Y(_03152_));
 sky130_fd_sc_hd__xnor2_2 _31549_ (.A(_03151_),
    .B(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__o21ba_2 _31550_ (.A1(_02746_),
    .A2(_02748_),
    .B1_N(_02745_),
    .X(_03154_));
 sky130_fd_sc_hd__xnor2_2 _31551_ (.A(_03153_),
    .B(_03154_),
    .Y(_03155_));
 sky130_fd_sc_hd__and2_2 _31552_ (.A(_03148_),
    .B(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__nor2_2 _31553_ (.A(_03148_),
    .B(_03155_),
    .Y(_03158_));
 sky130_fd_sc_hd__or2_2 _31554_ (.A(_03156_),
    .B(_03158_),
    .X(_03159_));
 sky130_fd_sc_hd__a21o_2 _31555_ (.A1(_02728_),
    .A2(_03142_),
    .B1(_03159_),
    .X(_03160_));
 sky130_fd_sc_hd__nand3_2 _31556_ (.A(_02728_),
    .B(_03142_),
    .C(_03159_),
    .Y(_03161_));
 sky130_fd_sc_hd__o211ai_2 _31557_ (.A1(_03141_),
    .A2(_02753_),
    .B1(_03160_),
    .C1(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__a211o_2 _31558_ (.A1(_03160_),
    .A2(_03161_),
    .B1(_03141_),
    .C1(_02753_),
    .X(_03163_));
 sky130_fd_sc_hd__and2_2 _31559_ (.A(_03162_),
    .B(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__xnor2_2 _31560_ (.A(_03140_),
    .B(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__nor2_2 _31561_ (.A(_02735_),
    .B(_02761_),
    .Y(_03166_));
 sky130_fd_sc_hd__or2_2 _31562_ (.A(_03165_),
    .B(_03166_),
    .X(_03167_));
 sky130_fd_sc_hd__nand2_2 _31563_ (.A(_03165_),
    .B(_03166_),
    .Y(_03169_));
 sky130_fd_sc_hd__nand2_2 _31564_ (.A(_03167_),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__or2_2 _31565_ (.A(_02797_),
    .B(_02799_),
    .X(_03171_));
 sky130_fd_sc_hd__and4_2 _31566_ (.A(iX[43]),
    .B(iX[44]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_03172_));
 sky130_fd_sc_hd__a22oi_2 _31567_ (.A1(iX[44]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[43]),
    .Y(_03173_));
 sky130_fd_sc_hd__nor2_2 _31568_ (.A(_03172_),
    .B(_03173_),
    .Y(_03174_));
 sky130_fd_sc_hd__nand2_2 _31569_ (.A(iX[42]),
    .B(iY[55]),
    .Y(_03175_));
 sky130_fd_sc_hd__xnor2_2 _31570_ (.A(_03174_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__and4_2 _31571_ (.A(iX[46]),
    .B(iX[47]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_03177_));
 sky130_fd_sc_hd__a22oi_2 _31572_ (.A1(iX[47]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[46]),
    .Y(_03178_));
 sky130_fd_sc_hd__nor2_2 _31573_ (.A(_03177_),
    .B(_03178_),
    .Y(_03180_));
 sky130_fd_sc_hd__nand2_2 _31574_ (.A(iX[45]),
    .B(iY[52]),
    .Y(_03181_));
 sky130_fd_sc_hd__xnor2_2 _31575_ (.A(_03180_),
    .B(_03181_),
    .Y(_03182_));
 sky130_fd_sc_hd__o21ba_2 _31576_ (.A1(_02773_),
    .A2(_02776_),
    .B1_N(_02772_),
    .X(_03183_));
 sky130_fd_sc_hd__xnor2_2 _31577_ (.A(_03182_),
    .B(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hd__and2_2 _31578_ (.A(_03176_),
    .B(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__nor2_2 _31579_ (.A(_03176_),
    .B(_03184_),
    .Y(_03186_));
 sky130_fd_sc_hd__or2_2 _31580_ (.A(_03185_),
    .B(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__or3_2 _31581_ (.A(_02784_),
    .B(_02789_),
    .C(_02790_),
    .X(_03188_));
 sky130_fd_sc_hd__o21ba_2 _31582_ (.A1(_02740_),
    .A2(_02743_),
    .B1_N(_02739_),
    .X(_03189_));
 sky130_fd_sc_hd__and4_2 _31583_ (.A(iY[47]),
    .B(iY[48]),
    .C(iX[49]),
    .D(iX[50]),
    .X(_03191_));
 sky130_fd_sc_hd__a22oi_2 _31584_ (.A1(iY[48]),
    .A2(iX[49]),
    .B1(iX[50]),
    .B2(iY[47]),
    .Y(_03192_));
 sky130_fd_sc_hd__nand2_2 _31585_ (.A(iX[48]),
    .B(iY[49]),
    .Y(_03193_));
 sky130_fd_sc_hd__o21a_2 _31586_ (.A1(_03191_),
    .A2(_03192_),
    .B1(_03193_),
    .X(_03194_));
 sky130_fd_sc_hd__nor3_2 _31587_ (.A(_03191_),
    .B(_03192_),
    .C(_03193_),
    .Y(_03195_));
 sky130_fd_sc_hd__nor2_2 _31588_ (.A(_03194_),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__xnor2_2 _31589_ (.A(_03189_),
    .B(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__o21ai_2 _31590_ (.A1(_02786_),
    .A2(_02790_),
    .B1(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__or3_2 _31591_ (.A(_02786_),
    .B(_02790_),
    .C(_03197_),
    .X(_03199_));
 sky130_fd_sc_hd__nand2_2 _31592_ (.A(_03198_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__a21oi_2 _31593_ (.A1(_03188_),
    .A2(_02793_),
    .B1(_03200_),
    .Y(_03202_));
 sky130_fd_sc_hd__and3_2 _31594_ (.A(_03188_),
    .B(_02793_),
    .C(_03200_),
    .X(_03203_));
 sky130_fd_sc_hd__or3_2 _31595_ (.A(_03187_),
    .B(_03202_),
    .C(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__o21ai_2 _31596_ (.A1(_03202_),
    .A2(_03203_),
    .B1(_03187_),
    .Y(_03205_));
 sky130_fd_sc_hd__nand2_2 _31597_ (.A(_03204_),
    .B(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__a21o_2 _31598_ (.A1(_02756_),
    .A2(_02758_),
    .B1(_03206_),
    .X(_03207_));
 sky130_fd_sc_hd__nand3_2 _31599_ (.A(_02756_),
    .B(_02758_),
    .C(_03206_),
    .Y(_03208_));
 sky130_fd_sc_hd__nand2_2 _31600_ (.A(_03207_),
    .B(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__xnor2_2 _31601_ (.A(_03171_),
    .B(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__xnor2_2 _31602_ (.A(_03170_),
    .B(_03210_),
    .Y(_03211_));
 sky130_fd_sc_hd__o21ai_2 _31603_ (.A1(_02764_),
    .A2(_02805_),
    .B1(_03211_),
    .Y(_03213_));
 sky130_fd_sc_hd__or3_2 _31604_ (.A(_02764_),
    .B(_02805_),
    .C(_03211_),
    .X(_03214_));
 sky130_fd_sc_hd__and2_2 _31605_ (.A(_03213_),
    .B(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__a21bo_2 _31606_ (.A1(_02830_),
    .A2(_02850_),
    .B1_N(_02849_),
    .X(_03216_));
 sky130_fd_sc_hd__or2b_2 _31607_ (.A(_02819_),
    .B_N(_02817_),
    .X(_03217_));
 sky130_fd_sc_hd__and4_2 _31608_ (.A(iX[37]),
    .B(iX[38]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_03218_));
 sky130_fd_sc_hd__a22oi_2 _31609_ (.A1(iX[38]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[37]),
    .Y(_03219_));
 sky130_fd_sc_hd__nor2_2 _31610_ (.A(_03218_),
    .B(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__nand2_2 _31611_ (.A(iX[36]),
    .B(iY[61]),
    .Y(_03221_));
 sky130_fd_sc_hd__xnor2_2 _31612_ (.A(_03220_),
    .B(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hd__o21ba_2 _31613_ (.A1(_02814_),
    .A2(_02816_),
    .B1_N(_02813_),
    .X(_03224_));
 sky130_fd_sc_hd__xnor2_2 _31614_ (.A(_03222_),
    .B(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__and2_2 _31615_ (.A(iX[35]),
    .B(iY[62]),
    .X(_03226_));
 sky130_fd_sc_hd__or2_2 _31616_ (.A(_03225_),
    .B(_03226_),
    .X(_03227_));
 sky130_fd_sc_hd__nand2_2 _31617_ (.A(_03225_),
    .B(_03226_),
    .Y(_03228_));
 sky130_fd_sc_hd__nand2_2 _31618_ (.A(_03227_),
    .B(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__a21oi_2 _31619_ (.A1(_03217_),
    .A2(_02823_),
    .B1(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__and3_2 _31620_ (.A(_03217_),
    .B(_02823_),
    .C(_03229_),
    .X(_03231_));
 sky130_fd_sc_hd__nor2_2 _31621_ (.A(_03230_),
    .B(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__nand2_2 _31622_ (.A(iX[34]),
    .B(iY[63]),
    .Y(_03233_));
 sky130_fd_sc_hd__xnor2_2 _31623_ (.A(_03232_),
    .B(_03233_),
    .Y(_03235_));
 sky130_fd_sc_hd__or2b_2 _31624_ (.A(_02835_),
    .B_N(_02841_),
    .X(_03236_));
 sky130_fd_sc_hd__or2b_2 _31625_ (.A(_02834_),
    .B_N(_02842_),
    .X(_03237_));
 sky130_fd_sc_hd__nand2_2 _31626_ (.A(_03236_),
    .B(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__and2b_2 _31627_ (.A_N(_02778_),
    .B(_02777_),
    .X(_03239_));
 sky130_fd_sc_hd__o21ba_2 _31628_ (.A1(_02837_),
    .A2(_02839_),
    .B1_N(_02836_),
    .X(_03240_));
 sky130_fd_sc_hd__o21ba_2 _31629_ (.A1(_02768_),
    .A2(_02770_),
    .B1_N(_02767_),
    .X(_03241_));
 sky130_fd_sc_hd__and4_2 _31630_ (.A(iX[40]),
    .B(iX[41]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_03242_));
 sky130_fd_sc_hd__a22oi_2 _31631_ (.A1(iX[41]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[40]),
    .Y(_03243_));
 sky130_fd_sc_hd__nor2_2 _31632_ (.A(_03242_),
    .B(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__nand2_2 _31633_ (.A(iX[39]),
    .B(iY[58]),
    .Y(_03246_));
 sky130_fd_sc_hd__xnor2_2 _31634_ (.A(_03244_),
    .B(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__xnor2_2 _31635_ (.A(_03241_),
    .B(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__xnor2_2 _31636_ (.A(_03240_),
    .B(_03248_),
    .Y(_03249_));
 sky130_fd_sc_hd__o21a_2 _31637_ (.A1(_03239_),
    .A2(_02780_),
    .B1(_03249_),
    .X(_03250_));
 sky130_fd_sc_hd__nor3_2 _31638_ (.A(_03239_),
    .B(_02780_),
    .C(_03249_),
    .Y(_03251_));
 sky130_fd_sc_hd__nor2_2 _31639_ (.A(_03250_),
    .B(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__xor2_2 _31640_ (.A(_03238_),
    .B(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__o21ai_2 _31641_ (.A1(_02844_),
    .A2(_02846_),
    .B1(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__or3_2 _31642_ (.A(_02844_),
    .B(_02846_),
    .C(_03253_),
    .X(_03255_));
 sky130_fd_sc_hd__and3_2 _31643_ (.A(_03235_),
    .B(_03254_),
    .C(_03255_),
    .X(_03257_));
 sky130_fd_sc_hd__a21oi_2 _31644_ (.A1(_03254_),
    .A2(_03255_),
    .B1(_03235_),
    .Y(_03258_));
 sky130_fd_sc_hd__nor2_2 _31645_ (.A(_03257_),
    .B(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__o21ai_2 _31646_ (.A1(_02801_),
    .A2(_02803_),
    .B1(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__or3_2 _31647_ (.A(_02801_),
    .B(_02803_),
    .C(_03259_),
    .X(_03261_));
 sky130_fd_sc_hd__and3_2 _31648_ (.A(_03216_),
    .B(_03260_),
    .C(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__a21oi_2 _31649_ (.A1(_03260_),
    .A2(_03261_),
    .B1(_03216_),
    .Y(_03263_));
 sky130_fd_sc_hd__nor2_2 _31650_ (.A(_03262_),
    .B(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__nand2_2 _31651_ (.A(_03215_),
    .B(_03264_),
    .Y(_03265_));
 sky130_fd_sc_hd__or2_2 _31652_ (.A(_03215_),
    .B(_03264_),
    .X(_03266_));
 sky130_fd_sc_hd__nand2_2 _31653_ (.A(_03265_),
    .B(_03266_),
    .Y(_03268_));
 sky130_fd_sc_hd__a21o_2 _31654_ (.A1(_02808_),
    .A2(_02860_),
    .B1(_03268_),
    .X(_03269_));
 sky130_fd_sc_hd__nand3_2 _31655_ (.A(_02808_),
    .B(_02860_),
    .C(_03268_),
    .Y(_03270_));
 sky130_fd_sc_hd__nand2_2 _31656_ (.A(_03269_),
    .B(_03270_),
    .Y(_03271_));
 sky130_fd_sc_hd__and2b_2 _31657_ (.A_N(_02858_),
    .B(_02811_),
    .X(_03272_));
 sky130_fd_sc_hd__nor2_2 _31658_ (.A(_02855_),
    .B(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__xnor2_2 _31659_ (.A(_03271_),
    .B(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__a21oi_2 _31660_ (.A1(_02866_),
    .A2(_02870_),
    .B1(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__and3_2 _31661_ (.A(_02866_),
    .B(_02870_),
    .C(_03274_),
    .X(_03276_));
 sky130_fd_sc_hd__or2_2 _31662_ (.A(_03275_),
    .B(_03276_),
    .X(_03277_));
 sky130_fd_sc_hd__o21ba_2 _31663_ (.A1(_02826_),
    .A2(_02828_),
    .B1_N(_02825_),
    .X(_03279_));
 sky130_fd_sc_hd__xnor2_2 _31664_ (.A(_03277_),
    .B(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__a21oi_2 _31665_ (.A1(_02875_),
    .A2(_02878_),
    .B1(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__nand3_2 _31666_ (.A(_02875_),
    .B(_02878_),
    .C(_03280_),
    .Y(_03282_));
 sky130_fd_sc_hd__or2b_2 _31667_ (.A(_03281_),
    .B_N(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__or2_2 _31668_ (.A(_02882_),
    .B(_02886_),
    .X(_03284_));
 sky130_fd_sc_hd__xnor2_2 _31669_ (.A(_03283_),
    .B(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hd__xnor2_2 _31670_ (.A(_03110_),
    .B(_03285_),
    .Y(_03286_));
 sky130_fd_sc_hd__xnor2_2 _31671_ (.A(_02912_),
    .B(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__and3_2 _31672_ (.A(_02911_),
    .B(_02890_),
    .C(_03287_),
    .X(_03288_));
 sky130_fd_sc_hd__a21o_2 _31673_ (.A1(_02911_),
    .A2(_02890_),
    .B1(_03287_),
    .X(_03290_));
 sky130_fd_sc_hd__and2b_2 _31674_ (.A_N(_03288_),
    .B(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__o21a_2 _31675_ (.A1(_02900_),
    .A2(_02903_),
    .B1(_02898_),
    .X(_03292_));
 sky130_fd_sc_hd__xnor2_2 _31676_ (.A(_03291_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__nand2_2 _31677_ (.A(_11590_),
    .B(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__nor2_2 _31678_ (.A(_11590_),
    .B(_03293_),
    .Y(_03295_));
 sky130_fd_sc_hd__inv_2 _31679_ (.A(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__nand2_2 _31680_ (.A(_03294_),
    .B(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__o21ai_2 _31681_ (.A1(_02908_),
    .A2(_02910_),
    .B1(_02905_),
    .Y(_03298_));
 sky130_fd_sc_hd__xnor2_2 _31682_ (.A(_03297_),
    .B(_03298_),
    .Y(oO[65]));
 sky130_fd_sc_hd__or2b_2 _31683_ (.A(_03285_),
    .B_N(_03110_),
    .X(_03300_));
 sky130_fd_sc_hd__nand2_2 _31684_ (.A(_02912_),
    .B(_03286_),
    .Y(_03301_));
 sky130_fd_sc_hd__and2_2 _31685_ (.A(_11777_),
    .B(_11778_),
    .X(_03302_));
 sky130_fd_sc_hd__nand2_2 _31686_ (.A(_02926_),
    .B(_02974_),
    .Y(_03303_));
 sky130_fd_sc_hd__or2b_2 _31687_ (.A(_02975_),
    .B_N(_02925_),
    .X(_03304_));
 sky130_fd_sc_hd__and2b_2 _31688_ (.A_N(_02947_),
    .B(_02950_),
    .X(_03305_));
 sky130_fd_sc_hd__a21oi_2 _31689_ (.A1(_02930_),
    .A2(_02951_),
    .B1(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__a21oi_2 _31690_ (.A1(_03303_),
    .A2(_03304_),
    .B1(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__and3_2 _31691_ (.A(_03303_),
    .B(_03304_),
    .C(_03306_),
    .X(_03308_));
 sky130_fd_sc_hd__nor2_2 _31692_ (.A(_03307_),
    .B(_03308_),
    .Y(_03309_));
 sky130_fd_sc_hd__or2b_2 _31693_ (.A(_02952_),
    .B_N(_02973_),
    .X(_03311_));
 sky130_fd_sc_hd__o21ai_2 _31694_ (.A1(_02969_),
    .A2(_02972_),
    .B1(_03311_),
    .Y(_03312_));
 sky130_fd_sc_hd__a21o_2 _31695_ (.A1(_02978_),
    .A2(_03019_),
    .B1(_03017_),
    .X(_03313_));
 sky130_fd_sc_hd__a21bo_2 _31696_ (.A1(_02932_),
    .A2(_02934_),
    .B1_N(_02931_),
    .X(_03314_));
 sky130_fd_sc_hd__or4b_2 _31697_ (.A(_16271_),
    .B(_18368_),
    .C(_02316_),
    .D_N(_01522_),
    .X(_03315_));
 sky130_fd_sc_hd__a2bb2o_2 _31698_ (.A1_N(_16271_),
    .A2_N(_02316_),
    .B1(_01522_),
    .B2(_18754_),
    .X(_03316_));
 sky130_fd_sc_hd__nand2_2 _31699_ (.A(_03315_),
    .B(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hd__buf_1 _31700_ (.A(_02322_),
    .X(_03318_));
 sky130_fd_sc_hd__nor2_2 _31701_ (.A(_18120_),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__xor2_2 _31702_ (.A(_03317_),
    .B(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__and4_2 _31703_ (.A(_02338_),
    .B(_01784_),
    .C(_00162_),
    .D(_00565_),
    .X(_03322_));
 sky130_fd_sc_hd__a22o_2 _31704_ (.A1(_01784_),
    .A2(_00162_),
    .B1(_00565_),
    .B2(_02338_),
    .X(_03323_));
 sky130_fd_sc_hd__or4b_2 _31705_ (.A(_00195_),
    .B(_00943_),
    .C(_03322_),
    .D_N(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__or4_2 _31706_ (.A(_00589_),
    .B(_00990_),
    .C(_02940_),
    .D(_02311_),
    .X(_03325_));
 sky130_fd_sc_hd__a22o_2 _31707_ (.A1(_01564_),
    .A2(_01733_),
    .B1(_03325_),
    .B2(_03323_),
    .X(_03326_));
 sky130_fd_sc_hd__buf_1 _31708_ (.A(_01510_),
    .X(_03327_));
 sky130_fd_sc_hd__a31o_2 _31709_ (.A1(_18754_),
    .A2(_03327_),
    .A3(_02937_),
    .B1(_02936_),
    .X(_03328_));
 sky130_fd_sc_hd__and3_2 _31710_ (.A(_03324_),
    .B(_03326_),
    .C(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__a21oi_2 _31711_ (.A1(_03324_),
    .A2(_03326_),
    .B1(_03328_),
    .Y(_03330_));
 sky130_fd_sc_hd__nor2_2 _31712_ (.A(_03329_),
    .B(_03330_),
    .Y(_03331_));
 sky130_fd_sc_hd__xor2_2 _31713_ (.A(_03320_),
    .B(_03331_),
    .X(_03333_));
 sky130_fd_sc_hd__o21bai_2 _31714_ (.A1(_02935_),
    .A2(_02945_),
    .B1_N(_02944_),
    .Y(_03334_));
 sky130_fd_sc_hd__xnor2_2 _31715_ (.A(_03333_),
    .B(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__xor2_2 _31716_ (.A(_03314_),
    .B(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__and2b_2 _31717_ (.A_N(_02965_),
    .B(_02959_),
    .X(_03337_));
 sky130_fd_sc_hd__a21o_2 _31718_ (.A1(_02958_),
    .A2(_02966_),
    .B1(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__and2b_2 _31719_ (.A_N(_02996_),
    .B(_02997_),
    .X(_03339_));
 sky130_fd_sc_hd__o21bai_2 _31720_ (.A1(_02988_),
    .A2(_02998_),
    .B1_N(_03339_),
    .Y(_03340_));
 sky130_fd_sc_hd__inv_2 _31721_ (.A(_18729_),
    .Y(_03341_));
 sky130_fd_sc_hd__or3b_2 _31722_ (.A(_00990_),
    .B(_03341_),
    .C_N(_02963_),
    .X(_03342_));
 sky130_fd_sc_hd__o21ai_2 _31723_ (.A1(_02961_),
    .A2(_02962_),
    .B1(_03342_),
    .Y(_03344_));
 sky130_fd_sc_hd__buf_1 _31724_ (.A(_18101_),
    .X(_03345_));
 sky130_fd_sc_hd__inv_2 _31725_ (.A(_02981_),
    .Y(_03346_));
 sky130_fd_sc_hd__a31o_2 _31726_ (.A1(_18157_),
    .A2(_03345_),
    .A3(_02986_),
    .B1(_03346_),
    .X(_03347_));
 sky130_fd_sc_hd__nand2_2 _31727_ (.A(_18157_),
    .B(_18732_),
    .Y(_03348_));
 sky130_fd_sc_hd__o32a_2 _31728_ (.A1(_15648_),
    .A2(_18111_),
    .A3(_18113_),
    .B1(_18343_),
    .B2(_01797_),
    .X(_03349_));
 sky130_fd_sc_hd__o21ba_2 _31729_ (.A1(_02962_),
    .A2(_03348_),
    .B1_N(_03349_),
    .X(_03350_));
 sky130_fd_sc_hd__nand2_2 _31730_ (.A(_01785_),
    .B(_02956_),
    .Y(_03351_));
 sky130_fd_sc_hd__xor2_2 _31731_ (.A(_03350_),
    .B(_03351_),
    .X(_03352_));
 sky130_fd_sc_hd__xnor2_2 _31732_ (.A(_03347_),
    .B(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__xnor2_2 _31733_ (.A(_03344_),
    .B(_03353_),
    .Y(_03355_));
 sky130_fd_sc_hd__xnor2_2 _31734_ (.A(_03340_),
    .B(_03355_),
    .Y(_03356_));
 sky130_fd_sc_hd__xor2_2 _31735_ (.A(_03338_),
    .B(_03356_),
    .X(_03357_));
 sky130_fd_sc_hd__and2b_2 _31736_ (.A_N(_02967_),
    .B(_02955_),
    .X(_03358_));
 sky130_fd_sc_hd__a21oi_2 _31737_ (.A1(_02954_),
    .A2(_02968_),
    .B1(_03358_),
    .Y(_03359_));
 sky130_fd_sc_hd__xnor2_2 _31738_ (.A(_03357_),
    .B(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__xnor2_2 _31739_ (.A(_03336_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__xor2_2 _31740_ (.A(_03313_),
    .B(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__xnor2_2 _31741_ (.A(_03312_),
    .B(_03362_),
    .Y(_03363_));
 sky130_fd_sc_hd__o21bai_2 _31742_ (.A1(_03011_),
    .A2(_03012_),
    .B1_N(_03014_),
    .Y(_03364_));
 sky130_fd_sc_hd__or2b_2 _31743_ (.A(_03022_),
    .B_N(_03041_),
    .X(_03366_));
 sky130_fd_sc_hd__or2b_2 _31744_ (.A(_03021_),
    .B_N(_03042_),
    .X(_03367_));
 sky130_fd_sc_hd__or4_2 _31745_ (.A(_02463_),
    .B(_02471_),
    .C(_18363_),
    .D(_17408_),
    .X(_03368_));
 sky130_fd_sc_hd__a22o_2 _31746_ (.A1(_02994_),
    .A2(_17394_),
    .B1(_02984_),
    .B2(_02983_),
    .X(_03369_));
 sky130_fd_sc_hd__and2_2 _31747_ (.A(_03368_),
    .B(_03369_),
    .X(_03370_));
 sky130_fd_sc_hd__nor2_2 _31748_ (.A(_01583_),
    .B(_17628_),
    .Y(_03371_));
 sky130_fd_sc_hd__xnor2_2 _31749_ (.A(_03370_),
    .B(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__nor2_2 _31750_ (.A(_15835_),
    .B(_01828_),
    .Y(_03373_));
 sky130_fd_sc_hd__and2_2 _31751_ (.A(_02990_),
    .B(_03373_),
    .X(_03374_));
 sky130_fd_sc_hd__nor2_2 _31752_ (.A(_02990_),
    .B(_03373_),
    .Y(_03375_));
 sky130_fd_sc_hd__nor2_2 _31753_ (.A(_03374_),
    .B(_03375_),
    .Y(_03377_));
 sky130_fd_sc_hd__buf_1 _31754_ (.A(_18181_),
    .X(_03378_));
 sky130_fd_sc_hd__nor2_2 _31755_ (.A(_03378_),
    .B(_16619_),
    .Y(_03379_));
 sky130_fd_sc_hd__xnor2_2 _31756_ (.A(_03377_),
    .B(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__or3b_2 _31757_ (.A(_03378_),
    .B(_01804_),
    .C_N(_02990_),
    .X(_03381_));
 sky130_fd_sc_hd__o21ai_2 _31758_ (.A1(_02991_),
    .A2(_02995_),
    .B1(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__and2b_2 _31759_ (.A_N(_03380_),
    .B(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__and2b_2 _31760_ (.A_N(_03382_),
    .B(_03380_),
    .X(_03384_));
 sky130_fd_sc_hd__nor2_2 _31761_ (.A(_03383_),
    .B(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__xnor2_2 _31762_ (.A(_03372_),
    .B(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__buf_1 _31763_ (.A(_15598_),
    .X(_03388_));
 sky130_fd_sc_hd__buf_1 _31764_ (.A(_01828_),
    .X(_03389_));
 sky130_fd_sc_hd__or3_2 _31765_ (.A(_03388_),
    .B(_03389_),
    .C(_03005_),
    .X(_03390_));
 sky130_fd_sc_hd__a21bo_2 _31766_ (.A1(_03002_),
    .A2(_03003_),
    .B1_N(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__or3b_2 _31767_ (.A(_15154_),
    .B(_01058_),
    .C_N(_03003_),
    .X(_03392_));
 sky130_fd_sc_hd__a22o_2 _31768_ (.A1(_15586_),
    .A2(_17488_),
    .B1(_17702_),
    .B2(_01033_),
    .X(_03393_));
 sky130_fd_sc_hd__nand2_2 _31769_ (.A(_03392_),
    .B(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__nor2_2 _31770_ (.A(_03388_),
    .B(_00255_),
    .Y(_03395_));
 sky130_fd_sc_hd__xnor2_2 _31771_ (.A(_03394_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__o21a_2 _31772_ (.A1(_03025_),
    .A2(_03030_),
    .B1(_03396_),
    .X(_03397_));
 sky130_fd_sc_hd__or3_2 _31773_ (.A(_03025_),
    .B(_03030_),
    .C(_03396_),
    .X(_03399_));
 sky130_fd_sc_hd__or2b_2 _31774_ (.A(_03397_),
    .B_N(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__xnor2_2 _31775_ (.A(_03391_),
    .B(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__a21oi_2 _31776_ (.A1(_03001_),
    .A2(_03007_),
    .B1(_03009_),
    .Y(_03402_));
 sky130_fd_sc_hd__xnor2_2 _31777_ (.A(_03401_),
    .B(_03402_),
    .Y(_03403_));
 sky130_fd_sc_hd__and2_2 _31778_ (.A(_03386_),
    .B(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__nor2_2 _31779_ (.A(_03386_),
    .B(_03403_),
    .Y(_03405_));
 sky130_fd_sc_hd__a211o_2 _31780_ (.A1(_03366_),
    .A2(_03367_),
    .B1(_03404_),
    .C1(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__o211ai_2 _31781_ (.A1(_03404_),
    .A2(_03405_),
    .B1(_03366_),
    .C1(_03367_),
    .Y(_03407_));
 sky130_fd_sc_hd__nand2_2 _31782_ (.A(_03406_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__xnor2_2 _31783_ (.A(_03364_),
    .B(_03408_),
    .Y(_03410_));
 sky130_fd_sc_hd__nor3_2 _31784_ (.A(_03029_),
    .B(_03030_),
    .C(_03040_),
    .Y(_03411_));
 sky130_fd_sc_hd__a21bo_2 _31785_ (.A1(_03044_),
    .A2(_03053_),
    .B1_N(_03052_),
    .X(_03412_));
 sky130_fd_sc_hd__nand2_2 _31786_ (.A(_03023_),
    .B(_18209_),
    .Y(_03413_));
 sky130_fd_sc_hd__nand2_2 _31787_ (.A(_14593_),
    .B(_18463_),
    .Y(_03414_));
 sky130_fd_sc_hd__or3_2 _31788_ (.A(_02608_),
    .B(_01066_),
    .C(_03414_),
    .X(_03415_));
 sky130_fd_sc_hd__o21ai_2 _31789_ (.A1(_02608_),
    .A2(_01066_),
    .B1(_03414_),
    .Y(_03416_));
 sky130_fd_sc_hd__nand2_2 _31790_ (.A(_03415_),
    .B(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__xor2_2 _31791_ (.A(_03413_),
    .B(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__nand2_2 _31792_ (.A(_13544_),
    .B(_00268_),
    .Y(_03419_));
 sky130_fd_sc_hd__nand2_2 _31793_ (.A(_17463_),
    .B(_02629_),
    .Y(_03421_));
 sky130_fd_sc_hd__xor2_2 _31794_ (.A(_03419_),
    .B(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__nand2_2 _31795_ (.A(_01647_),
    .B(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__a21o_2 _31796_ (.A1(_13889_),
    .A2(_01647_),
    .B1(_03422_),
    .X(_03424_));
 sky130_fd_sc_hd__o21ai_2 _31797_ (.A1(_02613_),
    .A2(_03423_),
    .B1(_03424_),
    .Y(_03425_));
 sky130_fd_sc_hd__o21ai_2 _31798_ (.A1(_03034_),
    .A2(_03035_),
    .B1(_03032_),
    .Y(_03426_));
 sky130_fd_sc_hd__xor2_2 _31799_ (.A(_03425_),
    .B(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__xor2_2 _31800_ (.A(_03418_),
    .B(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__xnor2_2 _31801_ (.A(_03412_),
    .B(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__o21a_2 _31802_ (.A1(_03038_),
    .A2(_03411_),
    .B1(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__nor3_2 _31803_ (.A(_03038_),
    .B(_03411_),
    .C(_03429_),
    .Y(_03432_));
 sky130_fd_sc_hd__nor2_2 _31804_ (.A(_03430_),
    .B(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__a31o_2 _31805_ (.A1(_02626_),
    .A2(_02629_),
    .A3(_03050_),
    .B1(_03047_),
    .X(_03434_));
 sky130_fd_sc_hd__nor2_2 _31806_ (.A(_02397_),
    .B(_02398_),
    .Y(_03435_));
 sky130_fd_sc_hd__and3_2 _31807_ (.A(_15677_),
    .B(_03435_),
    .C(_02644_),
    .X(_03436_));
 sky130_fd_sc_hd__a21o_2 _31808_ (.A1(_03057_),
    .A2(_03060_),
    .B1(_03436_),
    .X(_03437_));
 sky130_fd_sc_hd__buf_1 _31809_ (.A(_01650_),
    .X(_03438_));
 sky130_fd_sc_hd__nand2_2 _31810_ (.A(_02626_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__nor2_2 _31811_ (.A(_15646_),
    .B(_02391_),
    .Y(_03440_));
 sky130_fd_sc_hd__xnor2_2 _31812_ (.A(_03046_),
    .B(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__xor2_2 _31813_ (.A(_03439_),
    .B(_03441_),
    .X(_03443_));
 sky130_fd_sc_hd__xor2_2 _31814_ (.A(_03437_),
    .B(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__nand2_2 _31815_ (.A(_03434_),
    .B(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__or2_2 _31816_ (.A(_03434_),
    .B(_03444_),
    .X(_03446_));
 sky130_fd_sc_hd__and2_2 _31817_ (.A(_03445_),
    .B(_03446_),
    .X(_03447_));
 sky130_fd_sc_hd__o22a_2 _31818_ (.A1(_16625_),
    .A2(_03063_),
    .B1(_02663_),
    .B2(_11794_),
    .X(_03448_));
 sky130_fd_sc_hd__a21o_2 _31819_ (.A1(_12228_),
    .A2(_03064_),
    .B1(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__a21o_2 _31820_ (.A1(_11382_),
    .A2(_11586_),
    .B1(_03067_),
    .X(_03450_));
 sky130_fd_sc_hd__or2_2 _31821_ (.A(_03065_),
    .B(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__xnor2_2 _31822_ (.A(_03449_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__buf_1 _31823_ (.A(_03435_),
    .X(_03454_));
 sky130_fd_sc_hd__nand2_2 _31824_ (.A(_14649_),
    .B(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__and2_2 _31825_ (.A(_01880_),
    .B(_01881_),
    .X(_03456_));
 sky130_fd_sc_hd__buf_1 _31826_ (.A(_03456_),
    .X(_03457_));
 sky130_fd_sc_hd__buf_1 _31827_ (.A(_03457_),
    .X(_03458_));
 sky130_fd_sc_hd__nand2_2 _31828_ (.A(_00661_),
    .B(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__and3_2 _31829_ (.A(_00661_),
    .B(_03454_),
    .C(_02644_),
    .X(_03460_));
 sky130_fd_sc_hd__a21o_2 _31830_ (.A1(_03455_),
    .A2(_03459_),
    .B1(_03460_),
    .X(_03461_));
 sky130_fd_sc_hd__xor2_2 _31831_ (.A(_03452_),
    .B(_03461_),
    .X(_03462_));
 sky130_fd_sc_hd__nand2_2 _31832_ (.A(_02654_),
    .B(_02666_),
    .Y(_03463_));
 sky130_fd_sc_hd__o22ai_2 _31833_ (.A1(_03463_),
    .A2(_03066_),
    .B1(_03071_),
    .B2(_03062_),
    .Y(_03465_));
 sky130_fd_sc_hd__xor2_2 _31834_ (.A(_03462_),
    .B(_03465_),
    .X(_03466_));
 sky130_fd_sc_hd__xnor2_2 _31835_ (.A(_03447_),
    .B(_03466_),
    .Y(_03467_));
 sky130_fd_sc_hd__nor2_2 _31836_ (.A(_03072_),
    .B(_03075_),
    .Y(_03468_));
 sky130_fd_sc_hd__a21o_2 _31837_ (.A1(_03056_),
    .A2(_03076_),
    .B1(_03468_),
    .X(_03469_));
 sky130_fd_sc_hd__xnor2_2 _31838_ (.A(_03467_),
    .B(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__xnor2_2 _31839_ (.A(_03433_),
    .B(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__and2b_2 _31840_ (.A_N(_03080_),
    .B(_03077_),
    .X(_03472_));
 sky130_fd_sc_hd__a21oi_2 _31841_ (.A1(_03043_),
    .A2(_03082_),
    .B1(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__xor2_2 _31842_ (.A(_03471_),
    .B(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__xnor2_2 _31843_ (.A(_03410_),
    .B(_03474_),
    .Y(_03476_));
 sky130_fd_sc_hd__nor2_2 _31844_ (.A(_03083_),
    .B(_03085_),
    .Y(_03477_));
 sky130_fd_sc_hd__a21oi_2 _31845_ (.A1(_03020_),
    .A2(_03086_),
    .B1(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__xor2_2 _31846_ (.A(_03476_),
    .B(_03478_),
    .X(_03479_));
 sky130_fd_sc_hd__xnor2_2 _31847_ (.A(_03363_),
    .B(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__or2b_2 _31848_ (.A(_03089_),
    .B_N(_03087_),
    .X(_03481_));
 sky130_fd_sc_hd__o21ai_2 _31849_ (.A1(_02976_),
    .A2(_03090_),
    .B1(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__xnor2_2 _31850_ (.A(_03480_),
    .B(_03482_),
    .Y(_03483_));
 sky130_fd_sc_hd__xnor2_2 _31851_ (.A(_03309_),
    .B(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__nor2_2 _31852_ (.A(_03091_),
    .B(_03094_),
    .Y(_03485_));
 sky130_fd_sc_hd__a21oi_2 _31853_ (.A1(_02922_),
    .A2(_03095_),
    .B1(_03485_),
    .Y(_03487_));
 sky130_fd_sc_hd__xor2_2 _31854_ (.A(_03484_),
    .B(_03487_),
    .X(_03488_));
 sky130_fd_sc_hd__xnor2_2 _31855_ (.A(_02920_),
    .B(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__nor2_2 _31856_ (.A(_03096_),
    .B(_03098_),
    .Y(_03490_));
 sky130_fd_sc_hd__a21oi_2 _31857_ (.A1(_02514_),
    .A2(_03099_),
    .B1(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hd__xor2_2 _31858_ (.A(_03489_),
    .B(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__inv_2 _31859_ (.A(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__nor2_2 _31860_ (.A(_03101_),
    .B(_03102_),
    .Y(_03494_));
 sky130_fd_sc_hd__a21o_2 _31861_ (.A1(_02913_),
    .A2(_02914_),
    .B1(_03100_),
    .X(_03495_));
 sky130_fd_sc_hd__a21oi_2 _31862_ (.A1(_03107_),
    .A2(_03495_),
    .B1(_03102_),
    .Y(_03496_));
 sky130_fd_sc_hd__a41oi_2 _31863_ (.A1(_02691_),
    .A2(_03105_),
    .A3(_03106_),
    .A4(_03494_),
    .B1(_03496_),
    .Y(_03498_));
 sky130_fd_sc_hd__xnor2_2 _31864_ (.A(_03493_),
    .B(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hd__nor2_2 _31865_ (.A(_03277_),
    .B(_03279_),
    .Y(_03500_));
 sky130_fd_sc_hd__nand2_2 _31866_ (.A(_03140_),
    .B(_03164_),
    .Y(_03501_));
 sky130_fd_sc_hd__nor2_2 _31867_ (.A(_03119_),
    .B(_03121_),
    .Y(_03502_));
 sky130_fd_sc_hd__nand2_2 _31868_ (.A(iY[35]),
    .B(iX[63]),
    .Y(_03503_));
 sky130_fd_sc_hd__nor2_2 _31869_ (.A(_02704_),
    .B(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__a21oi_2 _31870_ (.A1(iY[37]),
    .A2(iX[61]),
    .B1(_01955_),
    .Y(_03505_));
 sky130_fd_sc_hd__and3_2 _31871_ (.A(iY[37]),
    .B(iX[62]),
    .C(_01373_),
    .X(_03506_));
 sky130_fd_sc_hd__nor2_2 _31872_ (.A(_03505_),
    .B(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__xnor2_2 _31873_ (.A(_03504_),
    .B(_03507_),
    .Y(_03509_));
 sky130_fd_sc_hd__a22oi_2 _31874_ (.A1(_03112_),
    .A2(_03113_),
    .B1(_03115_),
    .B2(_03118_),
    .Y(_03510_));
 sky130_fd_sc_hd__xnor2_2 _31875_ (.A(_03509_),
    .B(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__a31o_2 _31876_ (.A1(iY[40]),
    .A2(iX[57]),
    .A3(_03127_),
    .B1(_03126_),
    .X(_03512_));
 sky130_fd_sc_hd__nand2_2 _31877_ (.A(iY[38]),
    .B(iX[60]),
    .Y(_03513_));
 sky130_fd_sc_hd__nand2_2 _31878_ (.A(iY[39]),
    .B(iX[60]),
    .Y(_03514_));
 sky130_fd_sc_hd__nor2_2 _31879_ (.A(_03124_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__a21oi_2 _31880_ (.A1(_03125_),
    .A2(_03513_),
    .B1(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__nand2_2 _31881_ (.A(iY[40]),
    .B(iX[58]),
    .Y(_03517_));
 sky130_fd_sc_hd__xnor2_2 _31882_ (.A(_03516_),
    .B(_03517_),
    .Y(_03518_));
 sky130_fd_sc_hd__nand2_2 _31883_ (.A(_03117_),
    .B(_03518_),
    .Y(_03520_));
 sky130_fd_sc_hd__or2_2 _31884_ (.A(_03117_),
    .B(_03518_),
    .X(_03521_));
 sky130_fd_sc_hd__nand2_2 _31885_ (.A(_03520_),
    .B(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__xor2_2 _31886_ (.A(_03512_),
    .B(_03522_),
    .X(_03523_));
 sky130_fd_sc_hd__xor2_2 _31887_ (.A(_03511_),
    .B(_03523_),
    .X(_03524_));
 sky130_fd_sc_hd__o21a_2 _31888_ (.A1(_03502_),
    .A2(_03134_),
    .B1(_03524_),
    .X(_03525_));
 sky130_fd_sc_hd__nor3_2 _31889_ (.A(_03502_),
    .B(_03134_),
    .C(_03524_),
    .Y(_03526_));
 sky130_fd_sc_hd__nor2_2 _31890_ (.A(_03525_),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__and2b_2 _31891_ (.A_N(_03154_),
    .B(_03153_),
    .X(_03528_));
 sky130_fd_sc_hd__or2b_2 _31892_ (.A(_03132_),
    .B_N(_03123_),
    .X(_03529_));
 sky130_fd_sc_hd__and4_2 _31893_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[53]),
    .D(iX[54]),
    .X(_03531_));
 sky130_fd_sc_hd__a22oi_2 _31894_ (.A1(iY[45]),
    .A2(iX[53]),
    .B1(iX[54]),
    .B2(iY[44]),
    .Y(_03532_));
 sky130_fd_sc_hd__nor2_2 _31895_ (.A(_03531_),
    .B(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__nand2_2 _31896_ (.A(iY[46]),
    .B(iX[52]),
    .Y(_03534_));
 sky130_fd_sc_hd__xnor2_2 _31897_ (.A(_03533_),
    .B(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__and4_2 _31898_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[56]),
    .D(iX[57]),
    .X(_03536_));
 sky130_fd_sc_hd__a22oi_2 _31899_ (.A1(iY[42]),
    .A2(iX[56]),
    .B1(iX[57]),
    .B2(iY[41]),
    .Y(_03537_));
 sky130_fd_sc_hd__nor2_2 _31900_ (.A(_03536_),
    .B(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__nand2_2 _31901_ (.A(iY[43]),
    .B(iX[55]),
    .Y(_03539_));
 sky130_fd_sc_hd__xnor2_2 _31902_ (.A(_03538_),
    .B(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__o21ba_2 _31903_ (.A1(_03150_),
    .A2(_03152_),
    .B1_N(_03149_),
    .X(_03542_));
 sky130_fd_sc_hd__xnor2_2 _31904_ (.A(_03540_),
    .B(_03542_),
    .Y(_03543_));
 sky130_fd_sc_hd__xnor2_2 _31905_ (.A(_03535_),
    .B(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__a21o_2 _31906_ (.A1(_03130_),
    .A2(_03529_),
    .B1(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__nand3_2 _31907_ (.A(_03130_),
    .B(_03529_),
    .C(_03544_),
    .Y(_03546_));
 sky130_fd_sc_hd__o211ai_2 _31908_ (.A1(_03528_),
    .A2(_03156_),
    .B1(_03545_),
    .C1(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__a211o_2 _31909_ (.A1(_03545_),
    .A2(_03546_),
    .B1(_03528_),
    .C1(_03156_),
    .X(_03548_));
 sky130_fd_sc_hd__and2_2 _31910_ (.A(_03547_),
    .B(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__nor2_2 _31911_ (.A(_03527_),
    .B(_03549_),
    .Y(_03550_));
 sky130_fd_sc_hd__and2_2 _31912_ (.A(_03527_),
    .B(_03549_),
    .X(_03551_));
 sky130_fd_sc_hd__or2_2 _31913_ (.A(_03550_),
    .B(_03551_),
    .X(_03553_));
 sky130_fd_sc_hd__a21o_2 _31914_ (.A1(_03138_),
    .A2(_03501_),
    .B1(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__nand3_2 _31915_ (.A(_03138_),
    .B(_03501_),
    .C(_03553_),
    .Y(_03555_));
 sky130_fd_sc_hd__nand2_2 _31916_ (.A(_03554_),
    .B(_03555_),
    .Y(_03556_));
 sky130_fd_sc_hd__or2b_2 _31917_ (.A(_03202_),
    .B_N(_03204_),
    .X(_03557_));
 sky130_fd_sc_hd__and4_2 _31918_ (.A(iX[44]),
    .B(iX[45]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_03558_));
 sky130_fd_sc_hd__a22oi_2 _31919_ (.A1(iX[45]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[44]),
    .Y(_03559_));
 sky130_fd_sc_hd__nor2_2 _31920_ (.A(_03558_),
    .B(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__nand2_2 _31921_ (.A(iX[43]),
    .B(iY[55]),
    .Y(_03561_));
 sky130_fd_sc_hd__xnor2_2 _31922_ (.A(_03560_),
    .B(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__and4_2 _31923_ (.A(iX[47]),
    .B(iX[48]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_03564_));
 sky130_fd_sc_hd__a22oi_2 _31924_ (.A1(iX[48]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[47]),
    .Y(_03565_));
 sky130_fd_sc_hd__nor2_2 _31925_ (.A(_03564_),
    .B(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__nand2_2 _31926_ (.A(iX[46]),
    .B(iY[52]),
    .Y(_03567_));
 sky130_fd_sc_hd__xnor2_2 _31927_ (.A(_03566_),
    .B(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__o21ba_2 _31928_ (.A1(_03178_),
    .A2(_03181_),
    .B1_N(_03177_),
    .X(_03569_));
 sky130_fd_sc_hd__xnor2_2 _31929_ (.A(_03568_),
    .B(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__and2_2 _31930_ (.A(_03562_),
    .B(_03570_),
    .X(_03571_));
 sky130_fd_sc_hd__nor2_2 _31931_ (.A(_03562_),
    .B(_03570_),
    .Y(_03572_));
 sky130_fd_sc_hd__or2_2 _31932_ (.A(_03571_),
    .B(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__or3_2 _31933_ (.A(_03189_),
    .B(_03194_),
    .C(_03195_),
    .X(_03575_));
 sky130_fd_sc_hd__o21ba_2 _31934_ (.A1(_03144_),
    .A2(_03147_),
    .B1_N(_03143_),
    .X(_03576_));
 sky130_fd_sc_hd__and4_2 _31935_ (.A(iY[47]),
    .B(iY[48]),
    .C(iX[50]),
    .D(iX[51]),
    .X(_03577_));
 sky130_fd_sc_hd__a22oi_2 _31936_ (.A1(iY[48]),
    .A2(iX[50]),
    .B1(iX[51]),
    .B2(iY[47]),
    .Y(_03578_));
 sky130_fd_sc_hd__nand2_2 _31937_ (.A(iX[49]),
    .B(iY[49]),
    .Y(_03579_));
 sky130_fd_sc_hd__o21a_2 _31938_ (.A1(_03577_),
    .A2(_03578_),
    .B1(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__nor3_2 _31939_ (.A(_03577_),
    .B(_03578_),
    .C(_03579_),
    .Y(_03581_));
 sky130_fd_sc_hd__nor2_2 _31940_ (.A(_03580_),
    .B(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__xnor2_2 _31941_ (.A(_03576_),
    .B(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__o21ai_2 _31942_ (.A1(_03191_),
    .A2(_03195_),
    .B1(_03583_),
    .Y(_03584_));
 sky130_fd_sc_hd__or3_2 _31943_ (.A(_03191_),
    .B(_03195_),
    .C(_03583_),
    .X(_03586_));
 sky130_fd_sc_hd__nand2_2 _31944_ (.A(_03584_),
    .B(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__a21oi_2 _31945_ (.A1(_03575_),
    .A2(_03198_),
    .B1(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__and3_2 _31946_ (.A(_03575_),
    .B(_03198_),
    .C(_03587_),
    .X(_03589_));
 sky130_fd_sc_hd__or3_2 _31947_ (.A(_03573_),
    .B(_03588_),
    .C(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__o21ai_2 _31948_ (.A1(_03588_),
    .A2(_03589_),
    .B1(_03573_),
    .Y(_03591_));
 sky130_fd_sc_hd__nand2_2 _31949_ (.A(_03590_),
    .B(_03591_),
    .Y(_03592_));
 sky130_fd_sc_hd__a21oi_2 _31950_ (.A1(_03160_),
    .A2(_03162_),
    .B1(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__and3_2 _31951_ (.A(_03160_),
    .B(_03162_),
    .C(_03592_),
    .X(_03594_));
 sky130_fd_sc_hd__nor2_2 _31952_ (.A(_03593_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__xnor2_2 _31953_ (.A(_03557_),
    .B(_03595_),
    .Y(_03597_));
 sky130_fd_sc_hd__or2_2 _31954_ (.A(_03556_),
    .B(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__nand2_2 _31955_ (.A(_03556_),
    .B(_03597_),
    .Y(_03599_));
 sky130_fd_sc_hd__and2_2 _31956_ (.A(_03598_),
    .B(_03599_),
    .X(_03600_));
 sky130_fd_sc_hd__a21boi_2 _31957_ (.A1(_03169_),
    .A2(_03210_),
    .B1_N(_03167_),
    .Y(_03601_));
 sky130_fd_sc_hd__xnor2_2 _31958_ (.A(_03600_),
    .B(_03601_),
    .Y(_03602_));
 sky130_fd_sc_hd__a21boi_2 _31959_ (.A1(_03235_),
    .A2(_03255_),
    .B1_N(_03254_),
    .Y(_03603_));
 sky130_fd_sc_hd__or2b_2 _31960_ (.A(_03209_),
    .B_N(_03171_),
    .X(_03604_));
 sky130_fd_sc_hd__or2b_2 _31961_ (.A(_03224_),
    .B_N(_03222_),
    .X(_03605_));
 sky130_fd_sc_hd__and4_2 _31962_ (.A(iX[38]),
    .B(iX[39]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_03606_));
 sky130_fd_sc_hd__a22oi_2 _31963_ (.A1(iX[39]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[38]),
    .Y(_03608_));
 sky130_fd_sc_hd__nor2_2 _31964_ (.A(_03606_),
    .B(_03608_),
    .Y(_03609_));
 sky130_fd_sc_hd__nand2_2 _31965_ (.A(iX[37]),
    .B(iY[61]),
    .Y(_03610_));
 sky130_fd_sc_hd__xnor2_2 _31966_ (.A(_03609_),
    .B(_03610_),
    .Y(_03611_));
 sky130_fd_sc_hd__o21ba_2 _31967_ (.A1(_03219_),
    .A2(_03221_),
    .B1_N(_03218_),
    .X(_03612_));
 sky130_fd_sc_hd__xnor2_2 _31968_ (.A(_03611_),
    .B(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__and2_2 _31969_ (.A(iX[36]),
    .B(iY[62]),
    .X(_03614_));
 sky130_fd_sc_hd__or2_2 _31970_ (.A(_03613_),
    .B(_03614_),
    .X(_03615_));
 sky130_fd_sc_hd__nand2_2 _31971_ (.A(_03613_),
    .B(_03614_),
    .Y(_03616_));
 sky130_fd_sc_hd__nand2_2 _31972_ (.A(_03615_),
    .B(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__a21oi_2 _31973_ (.A1(_03605_),
    .A2(_03228_),
    .B1(_03617_),
    .Y(_03619_));
 sky130_fd_sc_hd__and3_2 _31974_ (.A(_03605_),
    .B(_03228_),
    .C(_03617_),
    .X(_03620_));
 sky130_fd_sc_hd__nor2_2 _31975_ (.A(_03619_),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__nand2_2 _31976_ (.A(iX[35]),
    .B(iY[63]),
    .Y(_03622_));
 sky130_fd_sc_hd__xnor2_2 _31977_ (.A(_03621_),
    .B(_03622_),
    .Y(_03623_));
 sky130_fd_sc_hd__or2b_2 _31978_ (.A(_03241_),
    .B_N(_03247_),
    .X(_03624_));
 sky130_fd_sc_hd__or2b_2 _31979_ (.A(_03240_),
    .B_N(_03248_),
    .X(_03625_));
 sky130_fd_sc_hd__and2b_2 _31980_ (.A_N(_03183_),
    .B(_03182_),
    .X(_03626_));
 sky130_fd_sc_hd__o21ba_2 _31981_ (.A1(_03243_),
    .A2(_03246_),
    .B1_N(_03242_),
    .X(_03627_));
 sky130_fd_sc_hd__o21ba_2 _31982_ (.A1(_03173_),
    .A2(_03175_),
    .B1_N(_03172_),
    .X(_03628_));
 sky130_fd_sc_hd__and4_2 _31983_ (.A(iX[41]),
    .B(iX[42]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_03630_));
 sky130_fd_sc_hd__a22oi_2 _31984_ (.A1(iX[42]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[41]),
    .Y(_03631_));
 sky130_fd_sc_hd__nor2_2 _31985_ (.A(_03630_),
    .B(_03631_),
    .Y(_03632_));
 sky130_fd_sc_hd__nand2_2 _31986_ (.A(iX[40]),
    .B(iY[58]),
    .Y(_03633_));
 sky130_fd_sc_hd__xnor2_2 _31987_ (.A(_03632_),
    .B(_03633_),
    .Y(_03634_));
 sky130_fd_sc_hd__xnor2_2 _31988_ (.A(_03628_),
    .B(_03634_),
    .Y(_03635_));
 sky130_fd_sc_hd__xnor2_2 _31989_ (.A(_03627_),
    .B(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__o21a_2 _31990_ (.A1(_03626_),
    .A2(_03185_),
    .B1(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__nor3_2 _31991_ (.A(_03626_),
    .B(_03185_),
    .C(_03636_),
    .Y(_03638_));
 sky130_fd_sc_hd__a211oi_2 _31992_ (.A1(_03624_),
    .A2(_03625_),
    .B1(_03637_),
    .C1(_03638_),
    .Y(_03639_));
 sky130_fd_sc_hd__o211a_2 _31993_ (.A1(_03637_),
    .A2(_03638_),
    .B1(_03624_),
    .C1(_03625_),
    .X(_03641_));
 sky130_fd_sc_hd__a21oi_2 _31994_ (.A1(_03238_),
    .A2(_03252_),
    .B1(_03250_),
    .Y(_03642_));
 sky130_fd_sc_hd__or3_2 _31995_ (.A(_03639_),
    .B(_03641_),
    .C(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__o21ai_2 _31996_ (.A1(_03639_),
    .A2(_03641_),
    .B1(_03642_),
    .Y(_03644_));
 sky130_fd_sc_hd__and3_2 _31997_ (.A(_03623_),
    .B(_03643_),
    .C(_03644_),
    .X(_03645_));
 sky130_fd_sc_hd__a21oi_2 _31998_ (.A1(_03643_),
    .A2(_03644_),
    .B1(_03623_),
    .Y(_03646_));
 sky130_fd_sc_hd__a211oi_2 _31999_ (.A1(_03207_),
    .A2(_03604_),
    .B1(_03645_),
    .C1(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__o211ai_2 _32000_ (.A1(_03645_),
    .A2(_03646_),
    .B1(_03207_),
    .C1(_03604_),
    .Y(_03648_));
 sky130_fd_sc_hd__or3b_2 _32001_ (.A(_03603_),
    .B(_03647_),
    .C_N(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__inv_2 _32002_ (.A(_03647_),
    .Y(_03650_));
 sky130_fd_sc_hd__a21bo_2 _32003_ (.A1(_03650_),
    .A2(_03648_),
    .B1_N(_03603_),
    .X(_03652_));
 sky130_fd_sc_hd__and2_2 _32004_ (.A(_03649_),
    .B(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__xnor2_2 _32005_ (.A(_03602_),
    .B(_03653_),
    .Y(_03654_));
 sky130_fd_sc_hd__a21oi_2 _32006_ (.A1(_03213_),
    .A2(_03265_),
    .B1(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__and3_2 _32007_ (.A(_03213_),
    .B(_03265_),
    .C(_03654_),
    .X(_03656_));
 sky130_fd_sc_hd__or2_2 _32008_ (.A(_03655_),
    .B(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__a21bo_2 _32009_ (.A1(_03216_),
    .A2(_03261_),
    .B1_N(_03260_),
    .X(_03658_));
 sky130_fd_sc_hd__xnor2_2 _32010_ (.A(_03657_),
    .B(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__o21ai_2 _32011_ (.A1(_03271_),
    .A2(_03273_),
    .B1(_03269_),
    .Y(_03660_));
 sky130_fd_sc_hd__xnor2_2 _32012_ (.A(_03659_),
    .B(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__a31o_2 _32013_ (.A1(iX[34]),
    .A2(iY[63]),
    .A3(_03232_),
    .B1(_03230_),
    .X(_03663_));
 sky130_fd_sc_hd__and2b_2 _32014_ (.A_N(_03661_),
    .B(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__and2b_2 _32015_ (.A_N(_03663_),
    .B(_03661_),
    .X(_03665_));
 sky130_fd_sc_hd__nor2_2 _32016_ (.A(_03664_),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__o21ai_2 _32017_ (.A1(_03275_),
    .A2(_03500_),
    .B1(_03666_),
    .Y(_03667_));
 sky130_fd_sc_hd__or3_2 _32018_ (.A(_03275_),
    .B(_03500_),
    .C(_03666_),
    .X(_03668_));
 sky130_fd_sc_hd__nand2_2 _32019_ (.A(_03667_),
    .B(_03668_),
    .Y(_03669_));
 sky130_fd_sc_hd__inv_2 _32020_ (.A(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__o31a_2 _32021_ (.A1(_02882_),
    .A2(_02886_),
    .A3(_03281_),
    .B1(_03282_),
    .X(_03671_));
 sky130_fd_sc_hd__xnor2_2 _32022_ (.A(_03670_),
    .B(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__xnor2_2 _32023_ (.A(_03499_),
    .B(_03672_),
    .Y(_03674_));
 sky130_fd_sc_hd__or2b_2 _32024_ (.A(_03302_),
    .B_N(_03674_),
    .X(_03675_));
 sky130_fd_sc_hd__or2b_2 _32025_ (.A(_03674_),
    .B_N(_03302_),
    .X(_03676_));
 sky130_fd_sc_hd__nand2_2 _32026_ (.A(_03675_),
    .B(_03676_),
    .Y(_03677_));
 sky130_fd_sc_hd__and3_2 _32027_ (.A(_03300_),
    .B(_03301_),
    .C(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__a21oi_2 _32028_ (.A1(_03300_),
    .A2(_03301_),
    .B1(_03677_),
    .Y(_03679_));
 sky130_fd_sc_hd__or2_2 _32029_ (.A(_03678_),
    .B(_03679_),
    .X(_03680_));
 sky130_fd_sc_hd__or2b_2 _32030_ (.A(_02900_),
    .B_N(_03291_),
    .X(_03681_));
 sky130_fd_sc_hd__a21oi_2 _32031_ (.A1(_02901_),
    .A2(_02902_),
    .B1(_03681_),
    .Y(_03682_));
 sky130_fd_sc_hd__o31a_2 _32032_ (.A1(_02892_),
    .A2(_02897_),
    .A3(_03288_),
    .B1(_03290_),
    .X(_03683_));
 sky130_fd_sc_hd__and2b_2 _32033_ (.A_N(_03682_),
    .B(_03683_),
    .X(_03685_));
 sky130_fd_sc_hd__xor2_2 _32034_ (.A(_03680_),
    .B(_03685_),
    .X(_03686_));
 sky130_fd_sc_hd__xor2_2 _32035_ (.A(_11808_),
    .B(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__nor2_2 _32036_ (.A(_02908_),
    .B(_03297_),
    .Y(_03688_));
 sky130_fd_sc_hd__o21a_2 _32037_ (.A1(_02507_),
    .A2(_02909_),
    .B1(_03688_),
    .X(_03689_));
 sky130_fd_sc_hd__a21oi_2 _32038_ (.A1(_02905_),
    .A2(_03294_),
    .B1(_03295_),
    .Y(_03690_));
 sky130_fd_sc_hd__nor2_2 _32039_ (.A(_03689_),
    .B(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__xnor2_2 _32040_ (.A(_03687_),
    .B(_03691_),
    .Y(oO[66]));
 sky130_fd_sc_hd__o21ba_2 _32041_ (.A1(_03680_),
    .A2(_03685_),
    .B1_N(_03679_),
    .X(_03692_));
 sky130_fd_sc_hd__xnor2_2 _32042_ (.A(_03669_),
    .B(_03671_),
    .Y(_03693_));
 sky130_fd_sc_hd__o21ai_2 _32043_ (.A1(_03499_),
    .A2(_03693_),
    .B1(_03675_),
    .Y(_03695_));
 sky130_fd_sc_hd__nand2_2 _32044_ (.A(_12038_),
    .B(_12039_),
    .Y(_03696_));
 sky130_fd_sc_hd__and2_2 _32045_ (.A(_03659_),
    .B(_03660_),
    .X(_03697_));
 sky130_fd_sc_hd__and2b_2 _32046_ (.A_N(_03657_),
    .B(_03658_),
    .X(_03698_));
 sky130_fd_sc_hd__a22oi_2 _32047_ (.A1(iY[37]),
    .A2(iX[62]),
    .B1(iX[63]),
    .B2(iY[36]),
    .Y(_03699_));
 sky130_fd_sc_hd__and3_2 _32048_ (.A(iY[37]),
    .B(iX[63]),
    .C(_01955_),
    .X(_03700_));
 sky130_fd_sc_hd__or2_2 _32049_ (.A(_03699_),
    .B(_03700_),
    .X(_03701_));
 sky130_fd_sc_hd__o21ba_2 _32050_ (.A1(_02704_),
    .A2(_03507_),
    .B1_N(_03503_),
    .X(_03702_));
 sky130_fd_sc_hd__or2b_2 _32051_ (.A(_03701_),
    .B_N(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__or2b_2 _32052_ (.A(_03702_),
    .B_N(_03701_),
    .X(_03704_));
 sky130_fd_sc_hd__nand2_2 _32053_ (.A(_03703_),
    .B(_03704_),
    .Y(_03706_));
 sky130_fd_sc_hd__a31o_2 _32054_ (.A1(iY[40]),
    .A2(iX[58]),
    .A3(_03516_),
    .B1(_03515_),
    .X(_03707_));
 sky130_fd_sc_hd__nand2_2 _32055_ (.A(iY[38]),
    .B(iX[61]),
    .Y(_03708_));
 sky130_fd_sc_hd__nand2_2 _32056_ (.A(iY[39]),
    .B(iX[61]),
    .Y(_03709_));
 sky130_fd_sc_hd__nor2_2 _32057_ (.A(_03513_),
    .B(_03709_),
    .Y(_03710_));
 sky130_fd_sc_hd__a21oi_2 _32058_ (.A1(_03514_),
    .A2(_03708_),
    .B1(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__nand2_2 _32059_ (.A(iY[40]),
    .B(iX[59]),
    .Y(_03712_));
 sky130_fd_sc_hd__xnor2_2 _32060_ (.A(_03711_),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__nand2_2 _32061_ (.A(_03506_),
    .B(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__or2_2 _32062_ (.A(_03506_),
    .B(_03713_),
    .X(_03715_));
 sky130_fd_sc_hd__nand2_2 _32063_ (.A(_03714_),
    .B(_03715_),
    .Y(_03717_));
 sky130_fd_sc_hd__xor2_2 _32064_ (.A(_03707_),
    .B(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__xnor2_2 _32065_ (.A(_03706_),
    .B(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__nor2_2 _32066_ (.A(_03511_),
    .B(_03523_),
    .Y(_03720_));
 sky130_fd_sc_hd__o21ba_2 _32067_ (.A1(_03509_),
    .A2(_03510_),
    .B1_N(_03720_),
    .X(_03721_));
 sky130_fd_sc_hd__xnor2_2 _32068_ (.A(_03719_),
    .B(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__and2b_2 _32069_ (.A_N(_03542_),
    .B(_03540_),
    .X(_03723_));
 sky130_fd_sc_hd__a21oi_2 _32070_ (.A1(_03535_),
    .A2(_03543_),
    .B1(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__or2b_2 _32071_ (.A(_03522_),
    .B_N(_03512_),
    .X(_03725_));
 sky130_fd_sc_hd__and4_2 _32072_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[54]),
    .D(iX[55]),
    .X(_03726_));
 sky130_fd_sc_hd__a22oi_2 _32073_ (.A1(iY[45]),
    .A2(iX[54]),
    .B1(iX[55]),
    .B2(iY[44]),
    .Y(_03728_));
 sky130_fd_sc_hd__nor2_2 _32074_ (.A(_03726_),
    .B(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__nand2_2 _32075_ (.A(iY[46]),
    .B(iX[53]),
    .Y(_03730_));
 sky130_fd_sc_hd__xnor2_2 _32076_ (.A(_03729_),
    .B(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__and4_2 _32077_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[57]),
    .D(iX[58]),
    .X(_03732_));
 sky130_fd_sc_hd__a22oi_2 _32078_ (.A1(iY[42]),
    .A2(iX[57]),
    .B1(iX[58]),
    .B2(iY[41]),
    .Y(_03733_));
 sky130_fd_sc_hd__nor2_2 _32079_ (.A(_03732_),
    .B(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand2_2 _32080_ (.A(iY[43]),
    .B(iX[56]),
    .Y(_03735_));
 sky130_fd_sc_hd__xnor2_2 _32081_ (.A(_03734_),
    .B(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__o21ba_2 _32082_ (.A1(_03537_),
    .A2(_03539_),
    .B1_N(_03536_),
    .X(_03737_));
 sky130_fd_sc_hd__xnor2_2 _32083_ (.A(_03736_),
    .B(_03737_),
    .Y(_03739_));
 sky130_fd_sc_hd__and2_2 _32084_ (.A(_03731_),
    .B(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__nor2_2 _32085_ (.A(_03731_),
    .B(_03739_),
    .Y(_03741_));
 sky130_fd_sc_hd__or2_2 _32086_ (.A(_03740_),
    .B(_03741_),
    .X(_03742_));
 sky130_fd_sc_hd__a21o_2 _32087_ (.A1(_03520_),
    .A2(_03725_),
    .B1(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__nand3_2 _32088_ (.A(_03520_),
    .B(_03725_),
    .C(_03742_),
    .Y(_03744_));
 sky130_fd_sc_hd__nand2_2 _32089_ (.A(_03743_),
    .B(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__xnor2_2 _32090_ (.A(_03724_),
    .B(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__and2_2 _32091_ (.A(_03722_),
    .B(_03746_),
    .X(_03747_));
 sky130_fd_sc_hd__nor2_2 _32092_ (.A(_03722_),
    .B(_03746_),
    .Y(_03748_));
 sky130_fd_sc_hd__nor2_2 _32093_ (.A(_03747_),
    .B(_03748_),
    .Y(_03750_));
 sky130_fd_sc_hd__o21a_2 _32094_ (.A1(_03525_),
    .A2(_03551_),
    .B1(_03750_),
    .X(_03751_));
 sky130_fd_sc_hd__nor3_2 _32095_ (.A(_03525_),
    .B(_03551_),
    .C(_03750_),
    .Y(_03752_));
 sky130_fd_sc_hd__nor2_2 _32096_ (.A(_03751_),
    .B(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__inv_2 _32097_ (.A(_03588_),
    .Y(_03754_));
 sky130_fd_sc_hd__and4_2 _32098_ (.A(iX[45]),
    .B(iX[46]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_03755_));
 sky130_fd_sc_hd__a22oi_2 _32099_ (.A1(iX[46]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[45]),
    .Y(_03756_));
 sky130_fd_sc_hd__nor2_2 _32100_ (.A(_03755_),
    .B(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__nand2_2 _32101_ (.A(iX[44]),
    .B(iY[55]),
    .Y(_03758_));
 sky130_fd_sc_hd__xnor2_2 _32102_ (.A(_03757_),
    .B(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__and4_2 _32103_ (.A(iX[48]),
    .B(iX[49]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_03761_));
 sky130_fd_sc_hd__a22oi_2 _32104_ (.A1(iX[49]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[48]),
    .Y(_03762_));
 sky130_fd_sc_hd__nor2_2 _32105_ (.A(_03761_),
    .B(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__nand2_2 _32106_ (.A(iX[47]),
    .B(iY[52]),
    .Y(_03764_));
 sky130_fd_sc_hd__xnor2_2 _32107_ (.A(_03763_),
    .B(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__o21ba_2 _32108_ (.A1(_03565_),
    .A2(_03567_),
    .B1_N(_03564_),
    .X(_03766_));
 sky130_fd_sc_hd__xnor2_2 _32109_ (.A(_03765_),
    .B(_03766_),
    .Y(_03767_));
 sky130_fd_sc_hd__and2_2 _32110_ (.A(_03759_),
    .B(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__nor2_2 _32111_ (.A(_03759_),
    .B(_03767_),
    .Y(_03769_));
 sky130_fd_sc_hd__or2_2 _32112_ (.A(_03768_),
    .B(_03769_),
    .X(_03770_));
 sky130_fd_sc_hd__or3_2 _32113_ (.A(_03576_),
    .B(_03580_),
    .C(_03581_),
    .X(_03772_));
 sky130_fd_sc_hd__o21ba_2 _32114_ (.A1(_03532_),
    .A2(_03534_),
    .B1_N(_03531_),
    .X(_03773_));
 sky130_fd_sc_hd__and4_2 _32115_ (.A(iY[47]),
    .B(iY[48]),
    .C(iX[51]),
    .D(iX[52]),
    .X(_03774_));
 sky130_fd_sc_hd__a22oi_2 _32116_ (.A1(iY[48]),
    .A2(iX[51]),
    .B1(iX[52]),
    .B2(iY[47]),
    .Y(_03775_));
 sky130_fd_sc_hd__nand2_2 _32117_ (.A(iY[49]),
    .B(iX[50]),
    .Y(_03776_));
 sky130_fd_sc_hd__o21a_2 _32118_ (.A1(_03774_),
    .A2(_03775_),
    .B1(_03776_),
    .X(_03777_));
 sky130_fd_sc_hd__nor3_2 _32119_ (.A(_03774_),
    .B(_03775_),
    .C(_03776_),
    .Y(_03778_));
 sky130_fd_sc_hd__nor2_2 _32120_ (.A(_03777_),
    .B(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hd__xnor2_2 _32121_ (.A(_03773_),
    .B(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__o21ai_2 _32122_ (.A1(_03577_),
    .A2(_03581_),
    .B1(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__or3_2 _32123_ (.A(_03577_),
    .B(_03581_),
    .C(_03780_),
    .X(_03783_));
 sky130_fd_sc_hd__nand2_2 _32124_ (.A(_03781_),
    .B(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__a21oi_2 _32125_ (.A1(_03772_),
    .A2(_03584_),
    .B1(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__and3_2 _32126_ (.A(_03772_),
    .B(_03584_),
    .C(_03784_),
    .X(_03786_));
 sky130_fd_sc_hd__or3_2 _32127_ (.A(_03770_),
    .B(_03785_),
    .C(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__o21ai_2 _32128_ (.A1(_03785_),
    .A2(_03786_),
    .B1(_03770_),
    .Y(_03788_));
 sky130_fd_sc_hd__nand2_2 _32129_ (.A(_03787_),
    .B(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__a21oi_2 _32130_ (.A1(_03545_),
    .A2(_03547_),
    .B1(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__and3_2 _32131_ (.A(_03545_),
    .B(_03547_),
    .C(_03789_),
    .X(_03791_));
 sky130_fd_sc_hd__a211oi_2 _32132_ (.A1(_03754_),
    .A2(_03590_),
    .B1(_03790_),
    .C1(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__o211a_2 _32133_ (.A1(_03790_),
    .A2(_03791_),
    .B1(_03754_),
    .C1(_03590_),
    .X(_03794_));
 sky130_fd_sc_hd__nor2_2 _32134_ (.A(_03792_),
    .B(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__and2_2 _32135_ (.A(_03753_),
    .B(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__nor2_2 _32136_ (.A(_03753_),
    .B(_03795_),
    .Y(_03797_));
 sky130_fd_sc_hd__or2_2 _32137_ (.A(_03796_),
    .B(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__a21o_2 _32138_ (.A1(_03554_),
    .A2(_03598_),
    .B1(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__nand3_2 _32139_ (.A(_03554_),
    .B(_03598_),
    .C(_03798_),
    .Y(_03800_));
 sky130_fd_sc_hd__nand2_2 _32140_ (.A(_03799_),
    .B(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__a21bo_2 _32141_ (.A1(_03623_),
    .A2(_03644_),
    .B1_N(_03643_),
    .X(_03802_));
 sky130_fd_sc_hd__and2_2 _32142_ (.A(_03557_),
    .B(_03595_),
    .X(_03803_));
 sky130_fd_sc_hd__or2b_2 _32143_ (.A(_03612_),
    .B_N(_03611_),
    .X(_03805_));
 sky130_fd_sc_hd__and4_2 _32144_ (.A(iX[39]),
    .B(iX[40]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_03806_));
 sky130_fd_sc_hd__a22oi_2 _32145_ (.A1(iX[40]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[39]),
    .Y(_03807_));
 sky130_fd_sc_hd__nor2_2 _32146_ (.A(_03806_),
    .B(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__nand2_2 _32147_ (.A(iX[38]),
    .B(iY[61]),
    .Y(_03809_));
 sky130_fd_sc_hd__xnor2_2 _32148_ (.A(_03808_),
    .B(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hd__o21ba_2 _32149_ (.A1(_03608_),
    .A2(_03610_),
    .B1_N(_03606_),
    .X(_03811_));
 sky130_fd_sc_hd__xnor2_2 _32150_ (.A(_03810_),
    .B(_03811_),
    .Y(_03812_));
 sky130_fd_sc_hd__and2_2 _32151_ (.A(iX[37]),
    .B(iY[62]),
    .X(_03813_));
 sky130_fd_sc_hd__nor2_2 _32152_ (.A(_03812_),
    .B(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__and2_2 _32153_ (.A(_03812_),
    .B(_03813_),
    .X(_03816_));
 sky130_fd_sc_hd__or2_2 _32154_ (.A(_03814_),
    .B(_03816_),
    .X(_03817_));
 sky130_fd_sc_hd__a21oi_2 _32155_ (.A1(_03805_),
    .A2(_03616_),
    .B1(_03817_),
    .Y(_03818_));
 sky130_fd_sc_hd__and3_2 _32156_ (.A(_03805_),
    .B(_03616_),
    .C(_03817_),
    .X(_03819_));
 sky130_fd_sc_hd__nor2_2 _32157_ (.A(_03818_),
    .B(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__nand2_2 _32158_ (.A(iX[36]),
    .B(iY[63]),
    .Y(_03821_));
 sky130_fd_sc_hd__xnor2_2 _32159_ (.A(_03820_),
    .B(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__or2b_2 _32160_ (.A(_03628_),
    .B_N(_03634_),
    .X(_03823_));
 sky130_fd_sc_hd__or2b_2 _32161_ (.A(_03627_),
    .B_N(_03635_),
    .X(_03824_));
 sky130_fd_sc_hd__and2b_2 _32162_ (.A_N(_03569_),
    .B(_03568_),
    .X(_03825_));
 sky130_fd_sc_hd__o21ba_2 _32163_ (.A1(_03631_),
    .A2(_03633_),
    .B1_N(_03630_),
    .X(_03827_));
 sky130_fd_sc_hd__o21ba_2 _32164_ (.A1(_03559_),
    .A2(_03561_),
    .B1_N(_03558_),
    .X(_03828_));
 sky130_fd_sc_hd__and4_2 _32165_ (.A(iX[42]),
    .B(iX[43]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_03829_));
 sky130_fd_sc_hd__a22oi_2 _32166_ (.A1(iX[43]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[42]),
    .Y(_03830_));
 sky130_fd_sc_hd__nor2_2 _32167_ (.A(_03829_),
    .B(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__nand2_2 _32168_ (.A(iX[41]),
    .B(iY[58]),
    .Y(_03832_));
 sky130_fd_sc_hd__xnor2_2 _32169_ (.A(_03831_),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__xnor2_2 _32170_ (.A(_03828_),
    .B(_03833_),
    .Y(_03834_));
 sky130_fd_sc_hd__xnor2_2 _32171_ (.A(_03827_),
    .B(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__o21a_2 _32172_ (.A1(_03825_),
    .A2(_03571_),
    .B1(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__nor3_2 _32173_ (.A(_03825_),
    .B(_03571_),
    .C(_03835_),
    .Y(_03838_));
 sky130_fd_sc_hd__a211oi_2 _32174_ (.A1(_03823_),
    .A2(_03824_),
    .B1(_03836_),
    .C1(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__o211a_2 _32175_ (.A1(_03836_),
    .A2(_03838_),
    .B1(_03823_),
    .C1(_03824_),
    .X(_03840_));
 sky130_fd_sc_hd__nor2_2 _32176_ (.A(_03637_),
    .B(_03639_),
    .Y(_03841_));
 sky130_fd_sc_hd__or3_2 _32177_ (.A(_03839_),
    .B(_03840_),
    .C(_03841_),
    .X(_03842_));
 sky130_fd_sc_hd__o21ai_2 _32178_ (.A1(_03839_),
    .A2(_03840_),
    .B1(_03841_),
    .Y(_03843_));
 sky130_fd_sc_hd__and3_2 _32179_ (.A(_03822_),
    .B(_03842_),
    .C(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__a21oi_2 _32180_ (.A1(_03842_),
    .A2(_03843_),
    .B1(_03822_),
    .Y(_03845_));
 sky130_fd_sc_hd__nor2_2 _32181_ (.A(_03844_),
    .B(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__o21a_2 _32182_ (.A1(_03593_),
    .A2(_03803_),
    .B1(_03846_),
    .X(_03847_));
 sky130_fd_sc_hd__nor3_2 _32183_ (.A(_03593_),
    .B(_03803_),
    .C(_03846_),
    .Y(_03849_));
 sky130_fd_sc_hd__or2_2 _32184_ (.A(_03847_),
    .B(_03849_),
    .X(_03850_));
 sky130_fd_sc_hd__xor2_2 _32185_ (.A(_03802_),
    .B(_03850_),
    .X(_03851_));
 sky130_fd_sc_hd__xor2_2 _32186_ (.A(_03801_),
    .B(_03851_),
    .X(_03852_));
 sky130_fd_sc_hd__and2b_2 _32187_ (.A_N(_03601_),
    .B(_03600_),
    .X(_03853_));
 sky130_fd_sc_hd__a21oi_2 _32188_ (.A1(_03602_),
    .A2(_03653_),
    .B1(_03853_),
    .Y(_03854_));
 sky130_fd_sc_hd__xnor2_2 _32189_ (.A(_03852_),
    .B(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__and2_2 _32190_ (.A(_03650_),
    .B(_03649_),
    .X(_03856_));
 sky130_fd_sc_hd__xnor2_2 _32191_ (.A(_03855_),
    .B(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__o21ai_2 _32192_ (.A1(_03655_),
    .A2(_03698_),
    .B1(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__or3_2 _32193_ (.A(_03655_),
    .B(_03698_),
    .C(_03857_),
    .X(_03860_));
 sky130_fd_sc_hd__nand2_2 _32194_ (.A(_03858_),
    .B(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__a31o_2 _32195_ (.A1(iX[35]),
    .A2(iY[63]),
    .A3(_03621_),
    .B1(_03619_),
    .X(_03862_));
 sky130_fd_sc_hd__xnor2_2 _32196_ (.A(_03861_),
    .B(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__o21ai_2 _32197_ (.A1(_03697_),
    .A2(_03664_),
    .B1(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__nor3_2 _32198_ (.A(_03697_),
    .B(_03664_),
    .C(_03863_),
    .Y(_03865_));
 sky130_fd_sc_hd__inv_2 _32199_ (.A(_03865_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand2_2 _32200_ (.A(_03864_),
    .B(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__a21bo_2 _32201_ (.A1(_03670_),
    .A2(_03671_),
    .B1_N(_03667_),
    .X(_03868_));
 sky130_fd_sc_hd__xor2_2 _32202_ (.A(_03867_),
    .B(_03868_),
    .X(_03869_));
 sky130_fd_sc_hd__nor2_2 _32203_ (.A(_03489_),
    .B(_03491_),
    .Y(_03871_));
 sky130_fd_sc_hd__o21bai_2 _32204_ (.A1(_03493_),
    .A2(_03498_),
    .B1_N(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__nor2_2 _32205_ (.A(_03484_),
    .B(_03487_),
    .Y(_03873_));
 sky130_fd_sc_hd__a21oi_2 _32206_ (.A1(_02920_),
    .A2(_03488_),
    .B1(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__or2b_2 _32207_ (.A(_03361_),
    .B_N(_03313_),
    .X(_03875_));
 sky130_fd_sc_hd__or2b_2 _32208_ (.A(_03362_),
    .B_N(_03312_),
    .X(_03876_));
 sky130_fd_sc_hd__and2b_2 _32209_ (.A_N(_03333_),
    .B(_03334_),
    .X(_03877_));
 sky130_fd_sc_hd__a21oi_2 _32210_ (.A1(_03314_),
    .A2(_03335_),
    .B1(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__a21oi_2 _32211_ (.A1(_03875_),
    .A2(_03876_),
    .B1(_03878_),
    .Y(_03879_));
 sky130_fd_sc_hd__and3_2 _32212_ (.A(_03875_),
    .B(_03876_),
    .C(_03878_),
    .X(_03880_));
 sky130_fd_sc_hd__nor2_2 _32213_ (.A(_03879_),
    .B(_03880_),
    .Y(_03882_));
 sky130_fd_sc_hd__and2b_2 _32214_ (.A_N(_03359_),
    .B(_03357_),
    .X(_03883_));
 sky130_fd_sc_hd__a21o_2 _32215_ (.A1(_03336_),
    .A2(_03360_),
    .B1(_03883_),
    .X(_03884_));
 sky130_fd_sc_hd__a21bo_2 _32216_ (.A1(_03364_),
    .A2(_03407_),
    .B1_N(_03406_),
    .X(_03885_));
 sky130_fd_sc_hd__a21bo_2 _32217_ (.A1(_03316_),
    .A2(_03319_),
    .B1_N(_03315_),
    .X(_03886_));
 sky130_fd_sc_hd__or4b_2 _32218_ (.A(_18368_),
    .B(_00195_),
    .C(_02316_),
    .D_N(_01521_),
    .X(_03887_));
 sky130_fd_sc_hd__a2bb2o_2 _32219_ (.A1_N(_18368_),
    .A2_N(_02316_),
    .B1(_01522_),
    .B2(_01564_),
    .X(_03888_));
 sky130_fd_sc_hd__nand2_2 _32220_ (.A(_03887_),
    .B(_03888_),
    .Y(_03889_));
 sky130_fd_sc_hd__nor2_2 _32221_ (.A(_16271_),
    .B(_02322_),
    .Y(_03890_));
 sky130_fd_sc_hd__xor2_2 _32222_ (.A(_03889_),
    .B(_03890_),
    .X(_03891_));
 sky130_fd_sc_hd__and4_2 _32223_ (.A(_01784_),
    .B(_01785_),
    .C(_00162_),
    .D(_00565_),
    .X(_03893_));
 sky130_fd_sc_hd__a22o_2 _32224_ (.A1(_01785_),
    .A2(_00162_),
    .B1(_00565_),
    .B2(_01784_),
    .X(_03894_));
 sky130_fd_sc_hd__or4b_2 _32225_ (.A(_00589_),
    .B(_00943_),
    .C(_03893_),
    .D_N(_03894_),
    .X(_03895_));
 sky130_fd_sc_hd__or4_2 _32226_ (.A(_00990_),
    .B(_16288_),
    .C(_02940_),
    .D(_01512_),
    .X(_03896_));
 sky130_fd_sc_hd__a22o_2 _32227_ (.A1(_02338_),
    .A2(_01733_),
    .B1(_03896_),
    .B2(_03894_),
    .X(_03897_));
 sky130_fd_sc_hd__a31o_2 _32228_ (.A1(_01564_),
    .A2(_01733_),
    .A3(_03323_),
    .B1(_03322_),
    .X(_03898_));
 sky130_fd_sc_hd__and3_2 _32229_ (.A(_03895_),
    .B(_03897_),
    .C(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__a21oi_2 _32230_ (.A1(_03895_),
    .A2(_03897_),
    .B1(_03898_),
    .Y(_03900_));
 sky130_fd_sc_hd__nor2_2 _32231_ (.A(_03899_),
    .B(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__xor2_2 _32232_ (.A(_03891_),
    .B(_03901_),
    .X(_03902_));
 sky130_fd_sc_hd__o21bai_2 _32233_ (.A1(_03320_),
    .A2(_03330_),
    .B1_N(_03329_),
    .Y(_03904_));
 sky130_fd_sc_hd__xnor2_2 _32234_ (.A(_03902_),
    .B(_03904_),
    .Y(_03905_));
 sky130_fd_sc_hd__xor2_2 _32235_ (.A(_03886_),
    .B(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__and2b_2 _32236_ (.A_N(_03352_),
    .B(_03347_),
    .X(_03907_));
 sky130_fd_sc_hd__a21o_2 _32237_ (.A1(_03344_),
    .A2(_03353_),
    .B1(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__o21ba_2 _32238_ (.A1(_03372_),
    .A2(_03384_),
    .B1_N(_03383_),
    .X(_03909_));
 sky130_fd_sc_hd__nor2_2 _32239_ (.A(_02962_),
    .B(_03348_),
    .Y(_03910_));
 sky130_fd_sc_hd__a31o_2 _32240_ (.A1(_01785_),
    .A2(_02956_),
    .A3(_03350_),
    .B1(_03910_),
    .X(_03911_));
 sky130_fd_sc_hd__a21bo_2 _32241_ (.A1(_03369_),
    .A2(_03371_),
    .B1_N(_03368_),
    .X(_03912_));
 sky130_fd_sc_hd__or3_2 _32242_ (.A(_01583_),
    .B(_18111_),
    .C(_18113_),
    .X(_03913_));
 sky130_fd_sc_hd__xor2_2 _32243_ (.A(_03348_),
    .B(_03913_),
    .X(_03915_));
 sky130_fd_sc_hd__nand2_2 _32244_ (.A(_00999_),
    .B(_18729_),
    .Y(_03916_));
 sky130_fd_sc_hd__xor2_2 _32245_ (.A(_03915_),
    .B(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__xnor2_2 _32246_ (.A(_03912_),
    .B(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__xnor2_2 _32247_ (.A(_03911_),
    .B(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__xnor2_2 _32248_ (.A(_03909_),
    .B(_03919_),
    .Y(_03920_));
 sky130_fd_sc_hd__xnor2_2 _32249_ (.A(_03908_),
    .B(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__and2b_2 _32250_ (.A_N(_03355_),
    .B(_03340_),
    .X(_03922_));
 sky130_fd_sc_hd__a21oi_2 _32251_ (.A1(_03338_),
    .A2(_03356_),
    .B1(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__xnor2_2 _32252_ (.A(_03921_),
    .B(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__xnor2_2 _32253_ (.A(_03906_),
    .B(_03924_),
    .Y(_03926_));
 sky130_fd_sc_hd__xor2_2 _32254_ (.A(_03885_),
    .B(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__xnor2_2 _32255_ (.A(_03884_),
    .B(_03927_),
    .Y(_03928_));
 sky130_fd_sc_hd__and2b_2 _32256_ (.A_N(_03402_),
    .B(_03401_),
    .X(_03929_));
 sky130_fd_sc_hd__or2_2 _32257_ (.A(_03929_),
    .B(_03404_),
    .X(_03930_));
 sky130_fd_sc_hd__and2b_2 _32258_ (.A_N(_03428_),
    .B(_03412_),
    .X(_03931_));
 sky130_fd_sc_hd__or4_2 _32259_ (.A(_02471_),
    .B(_18181_),
    .C(_18363_),
    .D(_17409_),
    .X(_03932_));
 sky130_fd_sc_hd__a22o_2 _32260_ (.A1(_02989_),
    .A2(_17394_),
    .B1(_02984_),
    .B2(_02994_),
    .X(_03933_));
 sky130_fd_sc_hd__and2_2 _32261_ (.A(_03932_),
    .B(_03933_),
    .X(_03934_));
 sky130_fd_sc_hd__nor2_2 _32262_ (.A(_02463_),
    .B(_17628_),
    .Y(_03935_));
 sky130_fd_sc_hd__xnor2_2 _32263_ (.A(_03934_),
    .B(_03935_),
    .Y(_03937_));
 sky130_fd_sc_hd__nor2_2 _32264_ (.A(_16257_),
    .B(_00255_),
    .Y(_03938_));
 sky130_fd_sc_hd__and2_2 _32265_ (.A(_03373_),
    .B(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__o22a_2 _32266_ (.A1(_01828_),
    .A2(_16258_),
    .B1(_00255_),
    .B2(_00996_),
    .X(_03940_));
 sky130_fd_sc_hd__nor2_2 _32267_ (.A(_03939_),
    .B(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__nor2_2 _32268_ (.A(_01832_),
    .B(_16619_),
    .Y(_03942_));
 sky130_fd_sc_hd__xnor2_2 _32269_ (.A(_03941_),
    .B(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__a21o_2 _32270_ (.A1(_03377_),
    .A2(_03379_),
    .B1(_03374_),
    .X(_03944_));
 sky130_fd_sc_hd__and2b_2 _32271_ (.A_N(_03943_),
    .B(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__and2b_2 _32272_ (.A_N(_03944_),
    .B(_03943_),
    .X(_03946_));
 sky130_fd_sc_hd__nor2_2 _32273_ (.A(_03945_),
    .B(_03946_),
    .Y(_03948_));
 sky130_fd_sc_hd__xnor2_2 _32274_ (.A(_03937_),
    .B(_03948_),
    .Y(_03949_));
 sky130_fd_sc_hd__a21bo_2 _32275_ (.A1(_03393_),
    .A2(_03395_),
    .B1_N(_03392_),
    .X(_03950_));
 sky130_fd_sc_hd__o21ai_2 _32276_ (.A1(_03413_),
    .A2(_03417_),
    .B1(_03415_),
    .Y(_03951_));
 sky130_fd_sc_hd__nor2_2 _32277_ (.A(_15173_),
    .B(_18200_),
    .Y(_03952_));
 sky130_fd_sc_hd__or3b_2 _32278_ (.A(_15155_),
    .B(_01058_),
    .C_N(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__a21o_2 _32279_ (.A1(_15586_),
    .A2(_17702_),
    .B1(_03952_),
    .X(_03954_));
 sky130_fd_sc_hd__nand2_2 _32280_ (.A(_03953_),
    .B(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__nor2_2 _32281_ (.A(_03388_),
    .B(_00649_),
    .Y(_03956_));
 sky130_fd_sc_hd__xor2_2 _32282_ (.A(_03955_),
    .B(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__xnor2_2 _32283_ (.A(_03951_),
    .B(_03957_),
    .Y(_03959_));
 sky130_fd_sc_hd__xnor2_2 _32284_ (.A(_03950_),
    .B(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__a21oi_2 _32285_ (.A1(_03391_),
    .A2(_03399_),
    .B1(_03397_),
    .Y(_03961_));
 sky130_fd_sc_hd__xor2_2 _32286_ (.A(_03960_),
    .B(_03961_),
    .X(_03962_));
 sky130_fd_sc_hd__xor2_2 _32287_ (.A(_03949_),
    .B(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__o21a_2 _32288_ (.A1(_03931_),
    .A2(_03430_),
    .B1(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__nor3_2 _32289_ (.A(_03931_),
    .B(_03430_),
    .C(_03963_),
    .Y(_03965_));
 sky130_fd_sc_hd__nor2_2 _32290_ (.A(_03964_),
    .B(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__xor2_2 _32291_ (.A(_03930_),
    .B(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__inv_2 _32292_ (.A(_03427_),
    .Y(_03968_));
 sky130_fd_sc_hd__or2b_2 _32293_ (.A(_03425_),
    .B_N(_03426_),
    .X(_03970_));
 sky130_fd_sc_hd__a21bo_2 _32294_ (.A1(_03418_),
    .A2(_03968_),
    .B1_N(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__nand2_2 _32295_ (.A(_03437_),
    .B(_03443_),
    .Y(_03972_));
 sky130_fd_sc_hd__buf_1 _32296_ (.A(_18463_),
    .X(_03973_));
 sky130_fd_sc_hd__nand2_2 _32297_ (.A(_03023_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__nor2_2 _32298_ (.A(_01605_),
    .B(_18211_),
    .Y(_03975_));
 sky130_fd_sc_hd__nand2_2 _32299_ (.A(_01039_),
    .B(_18460_),
    .Y(_03976_));
 sky130_fd_sc_hd__xnor2_2 _32300_ (.A(_03975_),
    .B(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__xnor2_2 _32301_ (.A(_03974_),
    .B(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__nand2_2 _32302_ (.A(_13889_),
    .B(_01862_),
    .Y(_03979_));
 sky130_fd_sc_hd__nand2_2 _32303_ (.A(_13544_),
    .B(_01650_),
    .Y(_03981_));
 sky130_fd_sc_hd__o22a_2 _32304_ (.A1(_18791_),
    .A2(_01070_),
    .B1(_01866_),
    .B2(_14626_),
    .X(_03982_));
 sky130_fd_sc_hd__o21ba_2 _32305_ (.A1(_03421_),
    .A2(_03981_),
    .B1_N(_03982_),
    .X(_03983_));
 sky130_fd_sc_hd__xnor2_2 _32306_ (.A(_03979_),
    .B(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__o22a_2 _32307_ (.A1(_03419_),
    .A2(_03421_),
    .B1(_03423_),
    .B2(_02613_),
    .X(_03985_));
 sky130_fd_sc_hd__xnor2_2 _32308_ (.A(_03984_),
    .B(_03985_),
    .Y(_03986_));
 sky130_fd_sc_hd__xnor2_2 _32309_ (.A(_03978_),
    .B(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__a21oi_2 _32310_ (.A1(_03972_),
    .A2(_03445_),
    .B1(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__nand3_2 _32311_ (.A(_03972_),
    .B(_03445_),
    .C(_03987_),
    .Y(_03989_));
 sky130_fd_sc_hd__or2b_2 _32312_ (.A(_03988_),
    .B_N(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__xnor2_2 _32313_ (.A(_03971_),
    .B(_03990_),
    .Y(_03992_));
 sky130_fd_sc_hd__o2bb2ai_2 _32314_ (.A1_N(_03046_),
    .A2_N(_03440_),
    .B1(_03441_),
    .B2(_03439_),
    .Y(_03993_));
 sky130_fd_sc_hd__buf_1 _32315_ (.A(_02641_),
    .X(_03994_));
 sky130_fd_sc_hd__and3_2 _32316_ (.A(_18192_),
    .B(_01880_),
    .C(_01881_),
    .X(_03995_));
 sky130_fd_sc_hd__a21oi_2 _32317_ (.A1(_14636_),
    .A2(_03994_),
    .B1(_03995_),
    .Y(_03996_));
 sky130_fd_sc_hd__a31o_2 _32318_ (.A1(_14636_),
    .A2(_03457_),
    .A3(_03440_),
    .B1(_03996_),
    .X(_03997_));
 sky130_fd_sc_hd__nor2_2 _32319_ (.A(_12852_),
    .B(_02647_),
    .Y(_03998_));
 sky130_fd_sc_hd__xnor2_2 _32320_ (.A(_03997_),
    .B(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hd__xor2_2 _32321_ (.A(_03460_),
    .B(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__xor2_2 _32322_ (.A(_03993_),
    .B(_04000_),
    .X(_04001_));
 sky130_fd_sc_hd__or2_2 _32323_ (.A(_03452_),
    .B(_03461_),
    .X(_04003_));
 sky130_fd_sc_hd__nand2_2 _32324_ (.A(_00661_),
    .B(_03454_),
    .Y(_04004_));
 sky130_fd_sc_hd__a31oi_2 _32325_ (.A1(_01877_),
    .A2(_01880_),
    .A3(_02394_),
    .B1(_02662_),
    .Y(_04005_));
 sky130_fd_sc_hd__a2bb2o_2 _32326_ (.A1_N(_18120_),
    .A2_N(_03063_),
    .B1(_04005_),
    .B2(_14649_),
    .X(_04006_));
 sky130_fd_sc_hd__o21ai_2 _32327_ (.A1(_12822_),
    .A2(_03068_),
    .B1(_04006_),
    .Y(_04007_));
 sky130_fd_sc_hd__or3_2 _32328_ (.A(_16625_),
    .B(_11794_),
    .C(_03067_),
    .X(_04008_));
 sky130_fd_sc_hd__o31ai_2 _32329_ (.A1(_03065_),
    .A2(_03448_),
    .A3(_03450_),
    .B1(_04008_),
    .Y(_04009_));
 sky130_fd_sc_hd__xor2_2 _32330_ (.A(_04007_),
    .B(_04009_),
    .X(_04010_));
 sky130_fd_sc_hd__xnor2_2 _32331_ (.A(_04004_),
    .B(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hd__xor2_2 _32332_ (.A(_04003_),
    .B(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__xnor2_2 _32333_ (.A(_04001_),
    .B(_04012_),
    .Y(_04014_));
 sky130_fd_sc_hd__nand2_2 _32334_ (.A(_03462_),
    .B(_03465_),
    .Y(_04015_));
 sky130_fd_sc_hd__a21bo_2 _32335_ (.A1(_03447_),
    .A2(_03466_),
    .B1_N(_04015_),
    .X(_04016_));
 sky130_fd_sc_hd__xnor2_2 _32336_ (.A(_04014_),
    .B(_04016_),
    .Y(_04017_));
 sky130_fd_sc_hd__xnor2_2 _32337_ (.A(_03992_),
    .B(_04017_),
    .Y(_04018_));
 sky130_fd_sc_hd__or2b_2 _32338_ (.A(_03467_),
    .B_N(_03469_),
    .X(_04019_));
 sky130_fd_sc_hd__a21bo_2 _32339_ (.A1(_03433_),
    .A2(_03470_),
    .B1_N(_04019_),
    .X(_04020_));
 sky130_fd_sc_hd__xnor2_2 _32340_ (.A(_04018_),
    .B(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__xnor2_2 _32341_ (.A(_03967_),
    .B(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__nor2_2 _32342_ (.A(_03471_),
    .B(_03473_),
    .Y(_04023_));
 sky130_fd_sc_hd__a21oi_2 _32343_ (.A1(_03410_),
    .A2(_03474_),
    .B1(_04023_),
    .Y(_04025_));
 sky130_fd_sc_hd__xor2_2 _32344_ (.A(_04022_),
    .B(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__xnor2_2 _32345_ (.A(_03928_),
    .B(_04026_),
    .Y(_04027_));
 sky130_fd_sc_hd__nor2_2 _32346_ (.A(_03476_),
    .B(_03478_),
    .Y(_04028_));
 sky130_fd_sc_hd__a21oi_2 _32347_ (.A1(_03363_),
    .A2(_03479_),
    .B1(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__xor2_2 _32348_ (.A(_04027_),
    .B(_04029_),
    .X(_04030_));
 sky130_fd_sc_hd__xnor2_2 _32349_ (.A(_03882_),
    .B(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__or2b_2 _32350_ (.A(_03480_),
    .B_N(_03482_),
    .X(_04032_));
 sky130_fd_sc_hd__a21boi_2 _32351_ (.A1(_03309_),
    .A2(_03483_),
    .B1_N(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__xor2_2 _32352_ (.A(_04031_),
    .B(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__xnor2_2 _32353_ (.A(_03307_),
    .B(_04034_),
    .Y(_04036_));
 sky130_fd_sc_hd__xor2_2 _32354_ (.A(_03874_),
    .B(_04036_),
    .X(_04037_));
 sky130_fd_sc_hd__xnor2_2 _32355_ (.A(_03872_),
    .B(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__and2b_2 _32356_ (.A_N(_03869_),
    .B(_04038_),
    .X(_04039_));
 sky130_fd_sc_hd__and2b_2 _32357_ (.A_N(_04038_),
    .B(_03869_),
    .X(_04040_));
 sky130_fd_sc_hd__nor2_2 _32358_ (.A(_04039_),
    .B(_04040_),
    .Y(_04041_));
 sky130_fd_sc_hd__xnor2_2 _32359_ (.A(_03696_),
    .B(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__xnor2_2 _32360_ (.A(_03695_),
    .B(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__xnor2_2 _32361_ (.A(_03692_),
    .B(_04043_),
    .Y(_04044_));
 sky130_fd_sc_hd__and2_2 _32362_ (.A(_11863_),
    .B(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__nor2_2 _32363_ (.A(_11863_),
    .B(_04044_),
    .Y(_04047_));
 sky130_fd_sc_hd__nor2_2 _32364_ (.A(_04045_),
    .B(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__nand2_2 _32365_ (.A(_11808_),
    .B(_03686_),
    .Y(_04049_));
 sky130_fd_sc_hd__o21ai_2 _32366_ (.A1(_03689_),
    .A2(_03690_),
    .B1(_03687_),
    .Y(_04050_));
 sky130_fd_sc_hd__nand2_2 _32367_ (.A(_04049_),
    .B(_04050_),
    .Y(_04051_));
 sky130_fd_sc_hd__xor2_2 _32368_ (.A(_04048_),
    .B(_04051_),
    .X(oO[67]));
 sky130_fd_sc_hd__inv_2 _32369_ (.A(_12211_),
    .Y(_04052_));
 sky130_fd_sc_hd__a21boi_2 _32370_ (.A1(_03874_),
    .A2(_04036_),
    .B1_N(_03871_),
    .Y(_04053_));
 sky130_fd_sc_hd__nor2_2 _32371_ (.A(_03874_),
    .B(_04036_),
    .Y(_04054_));
 sky130_fd_sc_hd__a311oi_2 _32372_ (.A1(_03492_),
    .A2(_03496_),
    .A3(_04037_),
    .B1(_04053_),
    .C1(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hd__nand2_2 _32373_ (.A(_03492_),
    .B(_04037_),
    .Y(_04057_));
 sky130_fd_sc_hd__inv_2 _32374_ (.A(_02691_),
    .Y(_04058_));
 sky130_fd_sc_hd__a2111o_2 _32375_ (.A1(_02693_),
    .A2(_02695_),
    .B1(_03104_),
    .C1(_04057_),
    .D1(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__or2b_2 _32376_ (.A(_03926_),
    .B_N(_03885_),
    .X(_04060_));
 sky130_fd_sc_hd__or2b_2 _32377_ (.A(_03927_),
    .B_N(_03884_),
    .X(_04061_));
 sky130_fd_sc_hd__and2b_2 _32378_ (.A_N(_03902_),
    .B(_03904_),
    .X(_04062_));
 sky130_fd_sc_hd__a21oi_2 _32379_ (.A1(_03886_),
    .A2(_03905_),
    .B1(_04062_),
    .Y(_04063_));
 sky130_fd_sc_hd__a21oi_2 _32380_ (.A1(_04060_),
    .A2(_04061_),
    .B1(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__and3_2 _32381_ (.A(_04060_),
    .B(_04061_),
    .C(_04063_),
    .X(_04065_));
 sky130_fd_sc_hd__nor2_2 _32382_ (.A(_04064_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__and2b_2 _32383_ (.A_N(_03923_),
    .B(_03921_),
    .X(_04068_));
 sky130_fd_sc_hd__a21o_2 _32384_ (.A1(_03906_),
    .A2(_03924_),
    .B1(_04068_),
    .X(_04069_));
 sky130_fd_sc_hd__a21o_2 _32385_ (.A1(_03930_),
    .A2(_03966_),
    .B1(_03964_),
    .X(_04070_));
 sky130_fd_sc_hd__a21bo_2 _32386_ (.A1(_03888_),
    .A2(_03890_),
    .B1_N(_03887_),
    .X(_04071_));
 sky130_fd_sc_hd__or4b_2 _32387_ (.A(_00195_),
    .B(_00589_),
    .C(_02316_),
    .D_N(_01521_),
    .X(_04072_));
 sky130_fd_sc_hd__a2bb2o_2 _32388_ (.A1_N(_00195_),
    .A2_N(_02316_),
    .B1(_01522_),
    .B2(_02338_),
    .X(_04073_));
 sky130_fd_sc_hd__nand2_2 _32389_ (.A(_04072_),
    .B(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__nor2_2 _32390_ (.A(_18368_),
    .B(_03318_),
    .Y(_04075_));
 sky130_fd_sc_hd__xor2_2 _32391_ (.A(_04074_),
    .B(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__or4_2 _32392_ (.A(_16288_),
    .B(_01797_),
    .C(_02940_),
    .D(_01512_),
    .X(_04077_));
 sky130_fd_sc_hd__a22o_2 _32393_ (.A1(_00999_),
    .A2(_00162_),
    .B1(_00565_),
    .B2(_01785_),
    .X(_04079_));
 sky130_fd_sc_hd__nand4_2 _32394_ (.A(_01784_),
    .B(_01733_),
    .C(_04077_),
    .D(_04079_),
    .Y(_04080_));
 sky130_fd_sc_hd__a22o_2 _32395_ (.A1(_01784_),
    .A2(_01733_),
    .B1(_04077_),
    .B2(_04079_),
    .X(_04081_));
 sky130_fd_sc_hd__a31o_2 _32396_ (.A1(_02338_),
    .A2(_01733_),
    .A3(_03894_),
    .B1(_03893_),
    .X(_04082_));
 sky130_fd_sc_hd__and3_2 _32397_ (.A(_04080_),
    .B(_04081_),
    .C(_04082_),
    .X(_04083_));
 sky130_fd_sc_hd__a21oi_2 _32398_ (.A1(_04080_),
    .A2(_04081_),
    .B1(_04082_),
    .Y(_04084_));
 sky130_fd_sc_hd__nor2_2 _32399_ (.A(_04083_),
    .B(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__xor2_2 _32400_ (.A(_04076_),
    .B(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__o21bai_2 _32401_ (.A1(_03891_),
    .A2(_03900_),
    .B1_N(_03899_),
    .Y(_04087_));
 sky130_fd_sc_hd__xnor2_2 _32402_ (.A(_04086_),
    .B(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__xor2_2 _32403_ (.A(_04071_),
    .B(_04088_),
    .X(_04090_));
 sky130_fd_sc_hd__and2b_2 _32404_ (.A_N(_03917_),
    .B(_03912_),
    .X(_04091_));
 sky130_fd_sc_hd__a21o_2 _32405_ (.A1(_03911_),
    .A2(_03918_),
    .B1(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__o21ba_2 _32406_ (.A1(_03937_),
    .A2(_03946_),
    .B1_N(_03945_),
    .X(_04093_));
 sky130_fd_sc_hd__nor2_2 _32407_ (.A(_03348_),
    .B(_03913_),
    .Y(_04094_));
 sky130_fd_sc_hd__a31o_2 _32408_ (.A1(_00999_),
    .A2(_02956_),
    .A3(_03915_),
    .B1(_04094_),
    .X(_04095_));
 sky130_fd_sc_hd__a21bo_2 _32409_ (.A1(_03933_),
    .A2(_03935_),
    .B1_N(_03932_),
    .X(_04096_));
 sky130_fd_sc_hd__nand2_2 _32410_ (.A(_02983_),
    .B(_18734_),
    .Y(_04097_));
 sky130_fd_sc_hd__o32ai_2 _32411_ (.A1(_02463_),
    .A2(_18111_),
    .A3(_18113_),
    .B1(_18343_),
    .B2(_01583_),
    .Y(_04098_));
 sky130_fd_sc_hd__o21a_2 _32412_ (.A1(_03913_),
    .A2(_04097_),
    .B1(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__nand2_2 _32413_ (.A(_18157_),
    .B(_02956_),
    .Y(_04101_));
 sky130_fd_sc_hd__xor2_2 _32414_ (.A(_04099_),
    .B(_04101_),
    .X(_04102_));
 sky130_fd_sc_hd__xnor2_2 _32415_ (.A(_04096_),
    .B(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__xnor2_2 _32416_ (.A(_04095_),
    .B(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__xnor2_2 _32417_ (.A(_04093_),
    .B(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__xnor2_2 _32418_ (.A(_04092_),
    .B(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__nand2_2 _32419_ (.A(_03909_),
    .B(_03919_),
    .Y(_04107_));
 sky130_fd_sc_hd__nor2_2 _32420_ (.A(_03909_),
    .B(_03919_),
    .Y(_04108_));
 sky130_fd_sc_hd__a21oi_2 _32421_ (.A1(_03908_),
    .A2(_04107_),
    .B1(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__xnor2_2 _32422_ (.A(_04106_),
    .B(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__xnor2_2 _32423_ (.A(_04090_),
    .B(_04110_),
    .Y(_04112_));
 sky130_fd_sc_hd__xor2_2 _32424_ (.A(_04070_),
    .B(_04112_),
    .X(_04113_));
 sky130_fd_sc_hd__xnor2_2 _32425_ (.A(_04069_),
    .B(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__nor2_2 _32426_ (.A(_03960_),
    .B(_03961_),
    .Y(_04115_));
 sky130_fd_sc_hd__a21oi_2 _32427_ (.A1(_03949_),
    .A2(_03962_),
    .B1(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__a21o_2 _32428_ (.A1(_03971_),
    .A2(_03989_),
    .B1(_03988_),
    .X(_04117_));
 sky130_fd_sc_hd__or2_2 _32429_ (.A(_16312_),
    .B(_16922_),
    .X(_04118_));
 sky130_fd_sc_hd__and3b_2 _32430_ (.A_N(_04118_),
    .B(_02984_),
    .C(_17460_),
    .X(_04119_));
 sky130_fd_sc_hd__o21a_2 _32431_ (.A1(_18181_),
    .A2(_17408_),
    .B1(_04118_),
    .X(_04120_));
 sky130_fd_sc_hd__nor2_2 _32432_ (.A(_04119_),
    .B(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__nor2_2 _32433_ (.A(_02471_),
    .B(_17628_),
    .Y(_04123_));
 sky130_fd_sc_hd__xnor2_2 _32434_ (.A(_04121_),
    .B(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__nor2_2 _32435_ (.A(_15835_),
    .B(_17007_),
    .Y(_04125_));
 sky130_fd_sc_hd__and2_2 _32436_ (.A(_03938_),
    .B(_04125_),
    .X(_04126_));
 sky130_fd_sc_hd__or2_2 _32437_ (.A(_03938_),
    .B(_04125_),
    .X(_04127_));
 sky130_fd_sc_hd__and2b_2 _32438_ (.A_N(_04126_),
    .B(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__nor2_2 _32439_ (.A(_01828_),
    .B(_16619_),
    .Y(_04129_));
 sky130_fd_sc_hd__xnor2_2 _32440_ (.A(_04128_),
    .B(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__a21o_2 _32441_ (.A1(_03941_),
    .A2(_03942_),
    .B1(_03939_),
    .X(_04131_));
 sky130_fd_sc_hd__and2b_2 _32442_ (.A_N(_04130_),
    .B(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__and2b_2 _32443_ (.A_N(_04131_),
    .B(_04130_),
    .X(_04134_));
 sky130_fd_sc_hd__nor2_2 _32444_ (.A(_04132_),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__xnor2_2 _32445_ (.A(_04124_),
    .B(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__a21bo_2 _32446_ (.A1(_03954_),
    .A2(_03956_),
    .B1_N(_03953_),
    .X(_04137_));
 sky130_fd_sc_hd__buf_1 _32447_ (.A(_01647_),
    .X(_04138_));
 sky130_fd_sc_hd__and3_2 _32448_ (.A(_14606_),
    .B(_18463_),
    .C(_03977_),
    .X(_04139_));
 sky130_fd_sc_hd__a31o_2 _32449_ (.A1(_01039_),
    .A2(_04138_),
    .A3(_03975_),
    .B1(_04139_),
    .X(_04140_));
 sky130_fd_sc_hd__nor2_2 _32450_ (.A(_15154_),
    .B(_18443_),
    .Y(_04141_));
 sky130_fd_sc_hd__o22a_2 _32451_ (.A1(_15154_),
    .A2(_18200_),
    .B1(_18443_),
    .B2(_15173_),
    .X(_04142_));
 sky130_fd_sc_hd__a21o_2 _32452_ (.A1(_03952_),
    .A2(_04141_),
    .B1(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__or2_2 _32453_ (.A(_03388_),
    .B(_01058_),
    .X(_04145_));
 sky130_fd_sc_hd__nand2_2 _32454_ (.A(_04143_),
    .B(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__or2_2 _32455_ (.A(_04143_),
    .B(_04145_),
    .X(_04147_));
 sky130_fd_sc_hd__nand2_2 _32456_ (.A(_04146_),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__xnor2_2 _32457_ (.A(_04140_),
    .B(_04148_),
    .Y(_04149_));
 sky130_fd_sc_hd__xnor2_2 _32458_ (.A(_04137_),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__and2b_2 _32459_ (.A_N(_03957_),
    .B(_03951_),
    .X(_04151_));
 sky130_fd_sc_hd__a21oi_2 _32460_ (.A1(_03950_),
    .A2(_03959_),
    .B1(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__xor2_2 _32461_ (.A(_04150_),
    .B(_04152_),
    .X(_04153_));
 sky130_fd_sc_hd__xor2_2 _32462_ (.A(_04136_),
    .B(_04153_),
    .X(_04154_));
 sky130_fd_sc_hd__xor2_2 _32463_ (.A(_04117_),
    .B(_04154_),
    .X(_04156_));
 sky130_fd_sc_hd__xnor2_2 _32464_ (.A(_04116_),
    .B(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__and2b_2 _32465_ (.A_N(_03985_),
    .B(_03984_),
    .X(_04158_));
 sky130_fd_sc_hd__a21oi_2 _32466_ (.A1(_03978_),
    .A2(_03986_),
    .B1(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__nand2_2 _32467_ (.A(_03460_),
    .B(_03999_),
    .Y(_04160_));
 sky130_fd_sc_hd__a21boi_2 _32468_ (.A1(_03993_),
    .A2(_04000_),
    .B1_N(_04160_),
    .Y(_04161_));
 sky130_fd_sc_hd__buf_1 _32469_ (.A(_00666_),
    .X(_04162_));
 sky130_fd_sc_hd__or3_2 _32470_ (.A(_01605_),
    .B(_04162_),
    .C(_03976_),
    .X(_04163_));
 sky130_fd_sc_hd__a22o_2 _32471_ (.A1(_14593_),
    .A2(_01647_),
    .B1(_00268_),
    .B2(_01039_),
    .X(_04164_));
 sky130_fd_sc_hd__nor2_2 _32472_ (.A(_01028_),
    .B(_01066_),
    .Y(_04165_));
 sky130_fd_sc_hd__a21o_2 _32473_ (.A1(_04163_),
    .A2(_04164_),
    .B1(_04165_),
    .X(_04167_));
 sky130_fd_sc_hd__nand3_2 _32474_ (.A(_04163_),
    .B(_04164_),
    .C(_04165_),
    .Y(_04168_));
 sky130_fd_sc_hd__nand2_2 _32475_ (.A(_04167_),
    .B(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__nor2_2 _32476_ (.A(_14641_),
    .B(_01087_),
    .Y(_04170_));
 sky130_fd_sc_hd__xnor2_2 _32477_ (.A(_03981_),
    .B(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__nor2_2 _32478_ (.A(_02613_),
    .B(_01070_),
    .Y(_04172_));
 sky130_fd_sc_hd__xnor2_2 _32479_ (.A(_04171_),
    .B(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__o22a_2 _32480_ (.A1(_03421_),
    .A2(_03981_),
    .B1(_03982_),
    .B2(_03979_),
    .X(_04174_));
 sky130_fd_sc_hd__xnor2_2 _32481_ (.A(_04173_),
    .B(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__xor2_2 _32482_ (.A(_04169_),
    .B(_04175_),
    .X(_04176_));
 sky130_fd_sc_hd__xnor2_2 _32483_ (.A(_04161_),
    .B(_04176_),
    .Y(_04178_));
 sky130_fd_sc_hd__xnor2_2 _32484_ (.A(_04159_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__or2_2 _32485_ (.A(_04004_),
    .B(_04010_),
    .X(_04180_));
 sky130_fd_sc_hd__buf_1 _32486_ (.A(_03063_),
    .X(_04181_));
 sky130_fd_sc_hd__a2bb2o_2 _32487_ (.A1_N(_16271_),
    .A2_N(_04181_),
    .B1(_04005_),
    .B2(_00661_),
    .X(_04182_));
 sky130_fd_sc_hd__o21a_2 _32488_ (.A1(_12823_),
    .A2(_03068_),
    .B1(_04182_),
    .X(_04183_));
 sky130_fd_sc_hd__a22o_2 _32489_ (.A1(_12755_),
    .A2(_03064_),
    .B1(_04006_),
    .B2(_04009_),
    .X(_04184_));
 sky130_fd_sc_hd__xnor2_2 _32490_ (.A(_04183_),
    .B(_04184_),
    .Y(_04185_));
 sky130_fd_sc_hd__xnor2_2 _32491_ (.A(_04180_),
    .B(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hd__buf_1 _32492_ (.A(_02647_),
    .X(_04187_));
 sky130_fd_sc_hd__nand2_2 _32493_ (.A(_14636_),
    .B(_03457_),
    .Y(_04189_));
 sky130_fd_sc_hd__or3_2 _32494_ (.A(_15646_),
    .B(_02391_),
    .C(_04189_),
    .X(_04190_));
 sky130_fd_sc_hd__o31ai_2 _32495_ (.A1(_12852_),
    .A2(_04187_),
    .A3(_03996_),
    .B1(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__nand2_2 _32496_ (.A(_02626_),
    .B(_03994_),
    .Y(_04192_));
 sky130_fd_sc_hd__and3_2 _32497_ (.A(_14636_),
    .B(_03435_),
    .C(_03995_),
    .X(_04193_));
 sky130_fd_sc_hd__o21a_2 _32498_ (.A1(_15646_),
    .A2(_02652_),
    .B1(_04189_),
    .X(_04194_));
 sky130_fd_sc_hd__nor2_2 _32499_ (.A(_04193_),
    .B(_04194_),
    .Y(_04195_));
 sky130_fd_sc_hd__xnor2_2 _32500_ (.A(_04192_),
    .B(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__nand2_2 _32501_ (.A(_04191_),
    .B(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__or2_2 _32502_ (.A(_04191_),
    .B(_04196_),
    .X(_04198_));
 sky130_fd_sc_hd__and2_2 _32503_ (.A(_04197_),
    .B(_04198_),
    .X(_04200_));
 sky130_fd_sc_hd__xnor2_2 _32504_ (.A(_04186_),
    .B(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__nor2_2 _32505_ (.A(_04003_),
    .B(_04011_),
    .Y(_04202_));
 sky130_fd_sc_hd__a21oi_2 _32506_ (.A1(_04001_),
    .A2(_04012_),
    .B1(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__xnor2_2 _32507_ (.A(_04201_),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__xnor2_2 _32508_ (.A(_04179_),
    .B(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__or2b_2 _32509_ (.A(_04014_),
    .B_N(_04016_),
    .X(_04206_));
 sky130_fd_sc_hd__a21bo_2 _32510_ (.A1(_03992_),
    .A2(_04017_),
    .B1_N(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__xnor2_2 _32511_ (.A(_04205_),
    .B(_04207_),
    .Y(_04208_));
 sky130_fd_sc_hd__xnor2_2 _32512_ (.A(_04157_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__or2b_2 _32513_ (.A(_04018_),
    .B_N(_04020_),
    .X(_04211_));
 sky130_fd_sc_hd__a21boi_2 _32514_ (.A1(_03967_),
    .A2(_04021_),
    .B1_N(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__xor2_2 _32515_ (.A(_04209_),
    .B(_04212_),
    .X(_04213_));
 sky130_fd_sc_hd__xnor2_2 _32516_ (.A(_04114_),
    .B(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__nor2_2 _32517_ (.A(_04022_),
    .B(_04025_),
    .Y(_04215_));
 sky130_fd_sc_hd__a21oi_2 _32518_ (.A1(_03928_),
    .A2(_04026_),
    .B1(_04215_),
    .Y(_04216_));
 sky130_fd_sc_hd__xor2_2 _32519_ (.A(_04214_),
    .B(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__xnor2_2 _32520_ (.A(_04066_),
    .B(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__nor2_2 _32521_ (.A(_04027_),
    .B(_04029_),
    .Y(_04219_));
 sky130_fd_sc_hd__a21oi_2 _32522_ (.A1(_03882_),
    .A2(_04030_),
    .B1(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__xor2_2 _32523_ (.A(_04218_),
    .B(_04220_),
    .X(_04222_));
 sky130_fd_sc_hd__xnor2_2 _32524_ (.A(_03879_),
    .B(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__nor2_2 _32525_ (.A(_04031_),
    .B(_04033_),
    .Y(_04224_));
 sky130_fd_sc_hd__a21oi_2 _32526_ (.A1(_03307_),
    .A2(_04034_),
    .B1(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__or2_2 _32527_ (.A(_04223_),
    .B(_04225_),
    .X(_04226_));
 sky130_fd_sc_hd__nand2_2 _32528_ (.A(_04223_),
    .B(_04225_),
    .Y(_04227_));
 sky130_fd_sc_hd__nand2_2 _32529_ (.A(_04226_),
    .B(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__a21o_2 _32530_ (.A1(_04055_),
    .A2(_04059_),
    .B1(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__nand3_2 _32531_ (.A(_04228_),
    .B(_04055_),
    .C(_04059_),
    .Y(_04230_));
 sky130_fd_sc_hd__nand2_2 _32532_ (.A(_04229_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__or2b_2 _32533_ (.A(_03861_),
    .B_N(_03862_),
    .X(_04233_));
 sky130_fd_sc_hd__or2b_2 _32534_ (.A(_03854_),
    .B_N(_03852_),
    .X(_04234_));
 sky130_fd_sc_hd__or2b_2 _32535_ (.A(_03856_),
    .B_N(_03855_),
    .X(_04235_));
 sky130_fd_sc_hd__nand2_2 _32536_ (.A(iY[37]),
    .B(iX[63]),
    .Y(_04236_));
 sky130_fd_sc_hd__a31o_2 _32537_ (.A1(iY[40]),
    .A2(iX[59]),
    .A3(_03711_),
    .B1(_03710_),
    .X(_04237_));
 sky130_fd_sc_hd__nand2_2 _32538_ (.A(iY[38]),
    .B(iX[62]),
    .Y(_04238_));
 sky130_fd_sc_hd__nand2_2 _32539_ (.A(iY[39]),
    .B(iX[62]),
    .Y(_04239_));
 sky130_fd_sc_hd__nor2_2 _32540_ (.A(_03708_),
    .B(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__a21oi_2 _32541_ (.A1(_03709_),
    .A2(_04238_),
    .B1(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__a21oi_2 _32542_ (.A1(iY[40]),
    .A2(iX[60]),
    .B1(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__and3_2 _32543_ (.A(iY[40]),
    .B(iX[60]),
    .C(_04241_),
    .X(_04244_));
 sky130_fd_sc_hd__nor2_2 _32544_ (.A(_04242_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__nand2_2 _32545_ (.A(_03700_),
    .B(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__or2_2 _32546_ (.A(_03700_),
    .B(_04245_),
    .X(_04247_));
 sky130_fd_sc_hd__nand2_2 _32547_ (.A(_04246_),
    .B(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__xor2_2 _32548_ (.A(_04237_),
    .B(_04248_),
    .X(_04249_));
 sky130_fd_sc_hd__or2_2 _32549_ (.A(_04236_),
    .B(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__nand2_2 _32550_ (.A(_04236_),
    .B(_04249_),
    .Y(_04251_));
 sky130_fd_sc_hd__nand2_2 _32551_ (.A(_04250_),
    .B(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__o21a_2 _32552_ (.A1(_03706_),
    .A2(_03718_),
    .B1(_03703_),
    .X(_04253_));
 sky130_fd_sc_hd__nor2_2 _32553_ (.A(_04252_),
    .B(_04253_),
    .Y(_04255_));
 sky130_fd_sc_hd__nand2_2 _32554_ (.A(_04252_),
    .B(_04253_),
    .Y(_04256_));
 sky130_fd_sc_hd__and2b_2 _32555_ (.A_N(_04255_),
    .B(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__and2b_2 _32556_ (.A_N(_03737_),
    .B(_03736_),
    .X(_04258_));
 sky130_fd_sc_hd__or2b_2 _32557_ (.A(_03717_),
    .B_N(_03707_),
    .X(_04259_));
 sky130_fd_sc_hd__and4_2 _32558_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[55]),
    .D(iX[56]),
    .X(_04260_));
 sky130_fd_sc_hd__a22oi_2 _32559_ (.A1(iY[45]),
    .A2(iX[55]),
    .B1(iX[56]),
    .B2(iY[44]),
    .Y(_04261_));
 sky130_fd_sc_hd__nor2_2 _32560_ (.A(_04260_),
    .B(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__nand2_2 _32561_ (.A(iY[46]),
    .B(iX[54]),
    .Y(_04263_));
 sky130_fd_sc_hd__xnor2_2 _32562_ (.A(_04262_),
    .B(_04263_),
    .Y(_04264_));
 sky130_fd_sc_hd__and4_2 _32563_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[58]),
    .D(iX[59]),
    .X(_04266_));
 sky130_fd_sc_hd__a22oi_2 _32564_ (.A1(iY[42]),
    .A2(iX[58]),
    .B1(iX[59]),
    .B2(iY[41]),
    .Y(_04267_));
 sky130_fd_sc_hd__nor2_2 _32565_ (.A(_04266_),
    .B(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__nand2_2 _32566_ (.A(iY[43]),
    .B(iX[57]),
    .Y(_04269_));
 sky130_fd_sc_hd__xnor2_2 _32567_ (.A(_04268_),
    .B(_04269_),
    .Y(_04270_));
 sky130_fd_sc_hd__o21ba_2 _32568_ (.A1(_03733_),
    .A2(_03735_),
    .B1_N(_03732_),
    .X(_04271_));
 sky130_fd_sc_hd__xnor2_2 _32569_ (.A(_04270_),
    .B(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__and2_2 _32570_ (.A(_04264_),
    .B(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__nor2_2 _32571_ (.A(_04264_),
    .B(_04272_),
    .Y(_04274_));
 sky130_fd_sc_hd__or2_2 _32572_ (.A(_04273_),
    .B(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__a21o_2 _32573_ (.A1(_03714_),
    .A2(_04259_),
    .B1(_04275_),
    .X(_04277_));
 sky130_fd_sc_hd__nand3_2 _32574_ (.A(_03714_),
    .B(_04259_),
    .C(_04275_),
    .Y(_04278_));
 sky130_fd_sc_hd__o211ai_2 _32575_ (.A1(_04258_),
    .A2(_03740_),
    .B1(_04277_),
    .C1(_04278_),
    .Y(_04279_));
 sky130_fd_sc_hd__a211o_2 _32576_ (.A1(_04277_),
    .A2(_04278_),
    .B1(_04258_),
    .C1(_03740_),
    .X(_04280_));
 sky130_fd_sc_hd__nand2_2 _32577_ (.A(_04279_),
    .B(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__xor2_2 _32578_ (.A(_04257_),
    .B(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__o21ba_2 _32579_ (.A1(_03719_),
    .A2(_03721_),
    .B1_N(_03748_),
    .X(_04283_));
 sky130_fd_sc_hd__xnor2_2 _32580_ (.A(_04282_),
    .B(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__or2b_2 _32581_ (.A(_03785_),
    .B_N(_03787_),
    .X(_04285_));
 sky130_fd_sc_hd__or2_2 _32582_ (.A(_03724_),
    .B(_03745_),
    .X(_04286_));
 sky130_fd_sc_hd__and4_2 _32583_ (.A(iX[46]),
    .B(iX[47]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_04288_));
 sky130_fd_sc_hd__a22oi_2 _32584_ (.A1(iX[47]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[46]),
    .Y(_04289_));
 sky130_fd_sc_hd__nor2_2 _32585_ (.A(_04288_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__nand2_2 _32586_ (.A(iX[45]),
    .B(iY[55]),
    .Y(_04291_));
 sky130_fd_sc_hd__xnor2_2 _32587_ (.A(_04290_),
    .B(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__and4_2 _32588_ (.A(iX[49]),
    .B(iX[50]),
    .C(iY[50]),
    .D(iY[51]),
    .X(_04293_));
 sky130_fd_sc_hd__a22oi_2 _32589_ (.A1(iX[50]),
    .A2(iY[50]),
    .B1(iY[51]),
    .B2(iX[49]),
    .Y(_04294_));
 sky130_fd_sc_hd__nor2_2 _32590_ (.A(_04293_),
    .B(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__nand2_2 _32591_ (.A(iX[48]),
    .B(iY[52]),
    .Y(_04296_));
 sky130_fd_sc_hd__xnor2_2 _32592_ (.A(_04295_),
    .B(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__o21ba_2 _32593_ (.A1(_03762_),
    .A2(_03764_),
    .B1_N(_03761_),
    .X(_04299_));
 sky130_fd_sc_hd__xnor2_2 _32594_ (.A(_04297_),
    .B(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__and2_2 _32595_ (.A(_04292_),
    .B(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__nor2_2 _32596_ (.A(_04292_),
    .B(_04300_),
    .Y(_04302_));
 sky130_fd_sc_hd__or2_2 _32597_ (.A(_04301_),
    .B(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__or3_2 _32598_ (.A(_03773_),
    .B(_03777_),
    .C(_03778_),
    .X(_04304_));
 sky130_fd_sc_hd__o21ba_2 _32599_ (.A1(_03728_),
    .A2(_03730_),
    .B1_N(_03726_),
    .X(_04305_));
 sky130_fd_sc_hd__and4_2 _32600_ (.A(iY[47]),
    .B(iY[48]),
    .C(iX[52]),
    .D(iX[53]),
    .X(_04306_));
 sky130_fd_sc_hd__a22oi_2 _32601_ (.A1(iY[48]),
    .A2(iX[52]),
    .B1(iX[53]),
    .B2(iY[47]),
    .Y(_04307_));
 sky130_fd_sc_hd__nand2_2 _32602_ (.A(iY[49]),
    .B(iX[51]),
    .Y(_04308_));
 sky130_fd_sc_hd__o21a_2 _32603_ (.A1(_04306_),
    .A2(_04307_),
    .B1(_04308_),
    .X(_04309_));
 sky130_fd_sc_hd__nor3_2 _32604_ (.A(_04306_),
    .B(_04307_),
    .C(_04308_),
    .Y(_04310_));
 sky130_fd_sc_hd__nor2_2 _32605_ (.A(_04309_),
    .B(_04310_),
    .Y(_04311_));
 sky130_fd_sc_hd__xnor2_2 _32606_ (.A(_04305_),
    .B(_04311_),
    .Y(_04312_));
 sky130_fd_sc_hd__o21ai_2 _32607_ (.A1(_03774_),
    .A2(_03778_),
    .B1(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__or3_2 _32608_ (.A(_03774_),
    .B(_03778_),
    .C(_04312_),
    .X(_04314_));
 sky130_fd_sc_hd__nand2_2 _32609_ (.A(_04313_),
    .B(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__a21oi_2 _32610_ (.A1(_04304_),
    .A2(_03781_),
    .B1(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__and3_2 _32611_ (.A(_04304_),
    .B(_03781_),
    .C(_04315_),
    .X(_04317_));
 sky130_fd_sc_hd__or3_2 _32612_ (.A(_04303_),
    .B(_04316_),
    .C(_04317_),
    .X(_04318_));
 sky130_fd_sc_hd__o21ai_2 _32613_ (.A1(_04316_),
    .A2(_04317_),
    .B1(_04303_),
    .Y(_04320_));
 sky130_fd_sc_hd__nand2_2 _32614_ (.A(_04318_),
    .B(_04320_),
    .Y(_04321_));
 sky130_fd_sc_hd__a21oi_2 _32615_ (.A1(_03743_),
    .A2(_04286_),
    .B1(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__and3_2 _32616_ (.A(_03743_),
    .B(_04286_),
    .C(_04321_),
    .X(_04323_));
 sky130_fd_sc_hd__nor2_2 _32617_ (.A(_04322_),
    .B(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__xnor2_2 _32618_ (.A(_04285_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__and2_2 _32619_ (.A(_04284_),
    .B(_04325_),
    .X(_04326_));
 sky130_fd_sc_hd__nor2_2 _32620_ (.A(_04284_),
    .B(_04325_),
    .Y(_04327_));
 sky130_fd_sc_hd__nor2_2 _32621_ (.A(_04326_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__o21ai_2 _32622_ (.A1(_03751_),
    .A2(_03796_),
    .B1(_04328_),
    .Y(_04329_));
 sky130_fd_sc_hd__or3_2 _32623_ (.A(_03751_),
    .B(_03796_),
    .C(_04328_),
    .X(_04331_));
 sky130_fd_sc_hd__and2_2 _32624_ (.A(_04329_),
    .B(_04331_),
    .X(_04332_));
 sky130_fd_sc_hd__a21boi_2 _32625_ (.A1(_03822_),
    .A2(_03843_),
    .B1_N(_03842_),
    .Y(_04333_));
 sky130_fd_sc_hd__and2b_2 _32626_ (.A_N(_03811_),
    .B(_03810_),
    .X(_04334_));
 sky130_fd_sc_hd__and4_2 _32627_ (.A(iX[40]),
    .B(iX[41]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_04335_));
 sky130_fd_sc_hd__a22oi_2 _32628_ (.A1(iX[41]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[40]),
    .Y(_04336_));
 sky130_fd_sc_hd__nor2_2 _32629_ (.A(_04335_),
    .B(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__nand2_2 _32630_ (.A(iX[39]),
    .B(iY[61]),
    .Y(_04338_));
 sky130_fd_sc_hd__xnor2_2 _32631_ (.A(_04337_),
    .B(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__o21ba_2 _32632_ (.A1(_03807_),
    .A2(_03809_),
    .B1_N(_03806_),
    .X(_04340_));
 sky130_fd_sc_hd__xnor2_2 _32633_ (.A(_04339_),
    .B(_04340_),
    .Y(_04342_));
 sky130_fd_sc_hd__and2_2 _32634_ (.A(iX[38]),
    .B(iY[62]),
    .X(_04343_));
 sky130_fd_sc_hd__or2_2 _32635_ (.A(_04342_),
    .B(_04343_),
    .X(_04344_));
 sky130_fd_sc_hd__nand2_2 _32636_ (.A(_04342_),
    .B(_04343_),
    .Y(_04345_));
 sky130_fd_sc_hd__o211a_2 _32637_ (.A1(_04334_),
    .A2(_03816_),
    .B1(_04344_),
    .C1(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_2 _32638_ (.A(_04344_),
    .B(_04345_),
    .Y(_04347_));
 sky130_fd_sc_hd__or3b_2 _32639_ (.A(_04334_),
    .B(_03816_),
    .C_N(_04347_),
    .X(_04348_));
 sky130_fd_sc_hd__and2b_2 _32640_ (.A_N(_04346_),
    .B(_04348_),
    .X(_04349_));
 sky130_fd_sc_hd__nand2_2 _32641_ (.A(iX[37]),
    .B(iY[63]),
    .Y(_04350_));
 sky130_fd_sc_hd__xnor2_2 _32642_ (.A(_04349_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__or2b_2 _32643_ (.A(_03828_),
    .B_N(_03833_),
    .X(_04353_));
 sky130_fd_sc_hd__or2b_2 _32644_ (.A(_03827_),
    .B_N(_03834_),
    .X(_04354_));
 sky130_fd_sc_hd__and2b_2 _32645_ (.A_N(_03766_),
    .B(_03765_),
    .X(_04355_));
 sky130_fd_sc_hd__o21ba_2 _32646_ (.A1(_03830_),
    .A2(_03832_),
    .B1_N(_03829_),
    .X(_04356_));
 sky130_fd_sc_hd__o21ba_2 _32647_ (.A1(_03756_),
    .A2(_03758_),
    .B1_N(_03755_),
    .X(_04357_));
 sky130_fd_sc_hd__and4_2 _32648_ (.A(iX[43]),
    .B(iX[44]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_04358_));
 sky130_fd_sc_hd__a22oi_2 _32649_ (.A1(iX[44]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[43]),
    .Y(_04359_));
 sky130_fd_sc_hd__nor2_2 _32650_ (.A(_04358_),
    .B(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__nand2_2 _32651_ (.A(iX[42]),
    .B(iY[58]),
    .Y(_04361_));
 sky130_fd_sc_hd__xnor2_2 _32652_ (.A(_04360_),
    .B(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__xnor2_2 _32653_ (.A(_04357_),
    .B(_04362_),
    .Y(_04364_));
 sky130_fd_sc_hd__xnor2_2 _32654_ (.A(_04356_),
    .B(_04364_),
    .Y(_04365_));
 sky130_fd_sc_hd__o21a_2 _32655_ (.A1(_04355_),
    .A2(_03768_),
    .B1(_04365_),
    .X(_04366_));
 sky130_fd_sc_hd__nor3_2 _32656_ (.A(_04355_),
    .B(_03768_),
    .C(_04365_),
    .Y(_04367_));
 sky130_fd_sc_hd__a211oi_2 _32657_ (.A1(_04353_),
    .A2(_04354_),
    .B1(_04366_),
    .C1(_04367_),
    .Y(_04368_));
 sky130_fd_sc_hd__o211a_2 _32658_ (.A1(_04366_),
    .A2(_04367_),
    .B1(_04353_),
    .C1(_04354_),
    .X(_04369_));
 sky130_fd_sc_hd__nor2_2 _32659_ (.A(_03836_),
    .B(_03839_),
    .Y(_04370_));
 sky130_fd_sc_hd__or3_2 _32660_ (.A(_04368_),
    .B(_04369_),
    .C(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__o21ai_2 _32661_ (.A1(_04368_),
    .A2(_04369_),
    .B1(_04370_),
    .Y(_04372_));
 sky130_fd_sc_hd__and3_2 _32662_ (.A(_04351_),
    .B(_04371_),
    .C(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__a21oi_2 _32663_ (.A1(_04371_),
    .A2(_04372_),
    .B1(_04351_),
    .Y(_04375_));
 sky130_fd_sc_hd__nor2_2 _32664_ (.A(_04373_),
    .B(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__o21a_2 _32665_ (.A1(_03790_),
    .A2(_03792_),
    .B1(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__nor3_2 _32666_ (.A(_03790_),
    .B(_03792_),
    .C(_04376_),
    .Y(_04378_));
 sky130_fd_sc_hd__nor2_2 _32667_ (.A(_04377_),
    .B(_04378_),
    .Y(_04379_));
 sky130_fd_sc_hd__xnor2_2 _32668_ (.A(_04333_),
    .B(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__nand2_2 _32669_ (.A(_04332_),
    .B(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__or2_2 _32670_ (.A(_04332_),
    .B(_04380_),
    .X(_04382_));
 sky130_fd_sc_hd__nand2_2 _32671_ (.A(_04381_),
    .B(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__o21a_2 _32672_ (.A1(_03801_),
    .A2(_03851_),
    .B1(_03799_),
    .X(_04384_));
 sky130_fd_sc_hd__or2_2 _32673_ (.A(_04383_),
    .B(_04384_),
    .X(_04386_));
 sky130_fd_sc_hd__nand2_2 _32674_ (.A(_04383_),
    .B(_04384_),
    .Y(_04387_));
 sky130_fd_sc_hd__nand2_2 _32675_ (.A(_04386_),
    .B(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__and2b_2 _32676_ (.A_N(_03850_),
    .B(_03802_),
    .X(_04389_));
 sky130_fd_sc_hd__nor2_2 _32677_ (.A(_03847_),
    .B(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__xnor2_2 _32678_ (.A(_04388_),
    .B(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hd__a21oi_2 _32679_ (.A1(_04234_),
    .A2(_04235_),
    .B1(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__and3_2 _32680_ (.A(_04234_),
    .B(_04235_),
    .C(_04391_),
    .X(_04393_));
 sky130_fd_sc_hd__or2_2 _32681_ (.A(_04392_),
    .B(_04393_),
    .X(_04394_));
 sky130_fd_sc_hd__a31o_2 _32682_ (.A1(iX[36]),
    .A2(iY[63]),
    .A3(_03820_),
    .B1(_03818_),
    .X(_04395_));
 sky130_fd_sc_hd__xor2_2 _32683_ (.A(_04394_),
    .B(_04395_),
    .X(_04397_));
 sky130_fd_sc_hd__a21o_2 _32684_ (.A1(_03858_),
    .A2(_04233_),
    .B1(_04397_),
    .X(_04398_));
 sky130_fd_sc_hd__nand3_2 _32685_ (.A(_03858_),
    .B(_04233_),
    .C(_04397_),
    .Y(_04399_));
 sky130_fd_sc_hd__nand2_2 _32686_ (.A(_04398_),
    .B(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__or2_2 _32687_ (.A(_03669_),
    .B(_03867_),
    .X(_04401_));
 sky130_fd_sc_hd__a2111o_2 _32688_ (.A1(_02699_),
    .A2(_02700_),
    .B1(_02885_),
    .C1(_03283_),
    .D1(_04401_),
    .X(_04402_));
 sky130_fd_sc_hd__o21ai_2 _32689_ (.A1(_02882_),
    .A2(_03281_),
    .B1(_03282_),
    .Y(_04403_));
 sky130_fd_sc_hd__o221a_2 _32690_ (.A1(_03667_),
    .A2(_03865_),
    .B1(_04401_),
    .B2(_04403_),
    .C1(_03864_),
    .X(_04404_));
 sky130_fd_sc_hd__nand2_2 _32691_ (.A(_04402_),
    .B(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__xnor2_2 _32692_ (.A(_04400_),
    .B(_04405_),
    .Y(_04406_));
 sky130_fd_sc_hd__nor2_2 _32693_ (.A(_04231_),
    .B(_04406_),
    .Y(_04408_));
 sky130_fd_sc_hd__and2_2 _32694_ (.A(_04231_),
    .B(_04406_),
    .X(_04409_));
 sky130_fd_sc_hd__nor2_2 _32695_ (.A(_04408_),
    .B(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__xnor2_2 _32696_ (.A(_04052_),
    .B(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__a21oi_2 _32697_ (.A1(_03696_),
    .A2(_04041_),
    .B1(_04040_),
    .Y(_04412_));
 sky130_fd_sc_hd__nor2_2 _32698_ (.A(_04411_),
    .B(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__and2_2 _32699_ (.A(_04411_),
    .B(_04412_),
    .X(_04414_));
 sky130_fd_sc_hd__or2_2 _32700_ (.A(_04413_),
    .B(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__and2b_2 _32701_ (.A_N(_03680_),
    .B(_04043_),
    .X(_04416_));
 sky130_fd_sc_hd__and2b_2 _32702_ (.A_N(_04042_),
    .B(_03695_),
    .X(_04417_));
 sky130_fd_sc_hd__nor2_2 _32703_ (.A(_03678_),
    .B(_03683_),
    .Y(_04419_));
 sky130_fd_sc_hd__or2b_2 _32704_ (.A(_03695_),
    .B_N(_04042_),
    .X(_04420_));
 sky130_fd_sc_hd__o31a_2 _32705_ (.A1(_03679_),
    .A2(_04417_),
    .A3(_04419_),
    .B1(_04420_),
    .X(_04421_));
 sky130_fd_sc_hd__a21oi_2 _32706_ (.A1(_03682_),
    .A2(_04416_),
    .B1(_04421_),
    .Y(_04422_));
 sky130_fd_sc_hd__xor2_2 _32707_ (.A(_04415_),
    .B(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__and2_2 _32708_ (.A(_12277_),
    .B(_04423_),
    .X(_04424_));
 sky130_fd_sc_hd__nor2_2 _32709_ (.A(_12277_),
    .B(_04423_),
    .Y(_04425_));
 sky130_fd_sc_hd__or2_2 _32710_ (.A(_04424_),
    .B(_04425_),
    .X(_04426_));
 sky130_fd_sc_hd__nand2_2 _32711_ (.A(_03687_),
    .B(_04048_),
    .Y(_04427_));
 sky130_fd_sc_hd__nand2_2 _32712_ (.A(_11863_),
    .B(_04044_),
    .Y(_04428_));
 sky130_fd_sc_hd__a21o_2 _32713_ (.A1(_04049_),
    .A2(_04428_),
    .B1(_04047_),
    .X(_04430_));
 sky130_fd_sc_hd__o21a_2 _32714_ (.A1(_03691_),
    .A2(_04427_),
    .B1(_04430_),
    .X(_04431_));
 sky130_fd_sc_hd__nor2_2 _32715_ (.A(_04426_),
    .B(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__and2_2 _32716_ (.A(_04426_),
    .B(_04431_),
    .X(_04433_));
 sky130_fd_sc_hd__nor2_2 _32717_ (.A(_04432_),
    .B(_04433_),
    .Y(oO[68]));
 sky130_fd_sc_hd__or2b_2 _32718_ (.A(_04112_),
    .B_N(_04070_),
    .X(_04434_));
 sky130_fd_sc_hd__or2b_2 _32719_ (.A(_04113_),
    .B_N(_04069_),
    .X(_04435_));
 sky130_fd_sc_hd__and2b_2 _32720_ (.A_N(_04086_),
    .B(_04087_),
    .X(_04436_));
 sky130_fd_sc_hd__a21oi_2 _32721_ (.A1(_04071_),
    .A2(_04088_),
    .B1(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__a21oi_2 _32722_ (.A1(_04434_),
    .A2(_04435_),
    .B1(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__and3_2 _32723_ (.A(_04434_),
    .B(_04435_),
    .C(_04437_),
    .X(_04440_));
 sky130_fd_sc_hd__nor2_2 _32724_ (.A(_04438_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__and2b_2 _32725_ (.A_N(_04109_),
    .B(_04106_),
    .X(_04442_));
 sky130_fd_sc_hd__a21o_2 _32726_ (.A1(_04090_),
    .A2(_04110_),
    .B1(_04442_),
    .X(_04443_));
 sky130_fd_sc_hd__or2b_2 _32727_ (.A(_04116_),
    .B_N(_04156_),
    .X(_04444_));
 sky130_fd_sc_hd__a21bo_2 _32728_ (.A1(_04117_),
    .A2(_04154_),
    .B1_N(_04444_),
    .X(_04445_));
 sky130_fd_sc_hd__a21bo_2 _32729_ (.A1(_04073_),
    .A2(_04075_),
    .B1_N(_04072_),
    .X(_04446_));
 sky130_fd_sc_hd__nor2_2 _32730_ (.A(_00589_),
    .B(_02316_),
    .Y(_04447_));
 sky130_fd_sc_hd__nand2_2 _32731_ (.A(_01784_),
    .B(_01522_),
    .Y(_04448_));
 sky130_fd_sc_hd__xnor2_2 _32732_ (.A(_04447_),
    .B(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__xor2_2 _32733_ (.A(_02320_),
    .B(_02321_),
    .X(_04451_));
 sky130_fd_sc_hd__nand2_2 _32734_ (.A(_01564_),
    .B(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__xnor2_2 _32735_ (.A(_04449_),
    .B(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__or4_2 _32736_ (.A(_01797_),
    .B(_01576_),
    .C(_02940_),
    .D(_01512_),
    .X(_04454_));
 sky130_fd_sc_hd__a22o_2 _32737_ (.A1(_18157_),
    .A2(_00162_),
    .B1(_00566_),
    .B2(_00999_),
    .X(_04455_));
 sky130_fd_sc_hd__nand2_2 _32738_ (.A(_04454_),
    .B(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hd__nand2_2 _32739_ (.A(_01785_),
    .B(_01733_),
    .Y(_04457_));
 sky130_fd_sc_hd__xnor2_2 _32740_ (.A(_04456_),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__and2_2 _32741_ (.A(_04077_),
    .B(_04080_),
    .X(_04459_));
 sky130_fd_sc_hd__xor2_2 _32742_ (.A(_04458_),
    .B(_04459_),
    .X(_04460_));
 sky130_fd_sc_hd__xnor2_2 _32743_ (.A(_04453_),
    .B(_04460_),
    .Y(_04462_));
 sky130_fd_sc_hd__o21bai_2 _32744_ (.A1(_04076_),
    .A2(_04084_),
    .B1_N(_04083_),
    .Y(_04463_));
 sky130_fd_sc_hd__xnor2_2 _32745_ (.A(_04462_),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__xor2_2 _32746_ (.A(_04446_),
    .B(_04464_),
    .X(_04465_));
 sky130_fd_sc_hd__or2b_2 _32747_ (.A(_04102_),
    .B_N(_04096_),
    .X(_04466_));
 sky130_fd_sc_hd__a21bo_2 _32748_ (.A1(_04095_),
    .A2(_04103_),
    .B1_N(_04466_),
    .X(_04467_));
 sky130_fd_sc_hd__o21bai_2 _32749_ (.A1(_04124_),
    .A2(_04134_),
    .B1_N(_04132_),
    .Y(_04468_));
 sky130_fd_sc_hd__buf_1 _32750_ (.A(_02956_),
    .X(_04469_));
 sky130_fd_sc_hd__nor2_2 _32751_ (.A(_03913_),
    .B(_04097_),
    .Y(_04470_));
 sky130_fd_sc_hd__a31o_2 _32752_ (.A1(_18157_),
    .A2(_04469_),
    .A3(_04098_),
    .B1(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__a31o_2 _32753_ (.A1(_02994_),
    .A2(_03345_),
    .A3(_04121_),
    .B1(_04119_),
    .X(_04473_));
 sky130_fd_sc_hd__or3_2 _32754_ (.A(_02471_),
    .B(_18111_),
    .C(_18113_),
    .X(_04474_));
 sky130_fd_sc_hd__xor2_2 _32755_ (.A(_04097_),
    .B(_04474_),
    .X(_04475_));
 sky130_fd_sc_hd__nand2_2 _32756_ (.A(_15888_),
    .B(_02956_),
    .Y(_04476_));
 sky130_fd_sc_hd__xnor2_2 _32757_ (.A(_04475_),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__xor2_2 _32758_ (.A(_04473_),
    .B(_04477_),
    .X(_04478_));
 sky130_fd_sc_hd__xnor2_2 _32759_ (.A(_04471_),
    .B(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__xor2_2 _32760_ (.A(_04468_),
    .B(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__xnor2_2 _32761_ (.A(_04467_),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__nand2_2 _32762_ (.A(_04093_),
    .B(_04104_),
    .Y(_04482_));
 sky130_fd_sc_hd__nor2_2 _32763_ (.A(_04093_),
    .B(_04104_),
    .Y(_04484_));
 sky130_fd_sc_hd__a21oi_2 _32764_ (.A1(_04092_),
    .A2(_04482_),
    .B1(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__xnor2_2 _32765_ (.A(_04481_),
    .B(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__xnor2_2 _32766_ (.A(_04465_),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__xor2_2 _32767_ (.A(_04445_),
    .B(_04487_),
    .X(_04488_));
 sky130_fd_sc_hd__xnor2_2 _32768_ (.A(_04443_),
    .B(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__nor2_2 _32769_ (.A(_04150_),
    .B(_04152_),
    .Y(_04490_));
 sky130_fd_sc_hd__a21o_2 _32770_ (.A1(_04136_),
    .A2(_04153_),
    .B1(_04490_),
    .X(_04491_));
 sky130_fd_sc_hd__and2b_2 _32771_ (.A_N(_04161_),
    .B(_04176_),
    .X(_04492_));
 sky130_fd_sc_hd__and2b_2 _32772_ (.A_N(_04159_),
    .B(_04178_),
    .X(_04493_));
 sky130_fd_sc_hd__or3_2 _32773_ (.A(_01828_),
    .B(_17409_),
    .C(_04118_),
    .X(_04495_));
 sky130_fd_sc_hd__a22o_2 _32774_ (.A1(_01040_),
    .A2(_17394_),
    .B1(_02984_),
    .B2(_00633_),
    .X(_04496_));
 sky130_fd_sc_hd__a22o_2 _32775_ (.A1(_02989_),
    .A2(_03345_),
    .B1(_04495_),
    .B2(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__nand4_2 _32776_ (.A(_02989_),
    .B(_03345_),
    .C(_04495_),
    .D(_04496_),
    .Y(_04498_));
 sky130_fd_sc_hd__nand2_2 _32777_ (.A(_04497_),
    .B(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__nor2_2 _32778_ (.A(_16258_),
    .B(_01058_),
    .Y(_04500_));
 sky130_fd_sc_hd__buf_1 _32779_ (.A(_01058_),
    .X(_04501_));
 sky130_fd_sc_hd__o22a_2 _32780_ (.A1(_16258_),
    .A2(_00649_),
    .B1(_04501_),
    .B2(_00996_),
    .X(_04502_));
 sky130_fd_sc_hd__a21oi_2 _32781_ (.A1(_04125_),
    .A2(_04500_),
    .B1(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__buf_1 _32782_ (.A(_00255_),
    .X(_04504_));
 sky130_fd_sc_hd__nor2_2 _32783_ (.A(_04504_),
    .B(_16619_),
    .Y(_04506_));
 sky130_fd_sc_hd__xnor2_2 _32784_ (.A(_04503_),
    .B(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__a21o_2 _32785_ (.A1(_04127_),
    .A2(_04129_),
    .B1(_04126_),
    .X(_04508_));
 sky130_fd_sc_hd__and2b_2 _32786_ (.A_N(_04507_),
    .B(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__and2b_2 _32787_ (.A_N(_04508_),
    .B(_04507_),
    .X(_04510_));
 sky130_fd_sc_hd__nor2_2 _32788_ (.A(_04509_),
    .B(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__xnor2_2 _32789_ (.A(_04499_),
    .B(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__a21bo_2 _32790_ (.A1(_03952_),
    .A2(_04141_),
    .B1_N(_04147_),
    .X(_04513_));
 sky130_fd_sc_hd__nor2_2 _32791_ (.A(_15173_),
    .B(_18211_),
    .Y(_04514_));
 sky130_fd_sc_hd__xor2_2 _32792_ (.A(_04141_),
    .B(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__nor2_2 _32793_ (.A(_03388_),
    .B(_18200_),
    .Y(_04517_));
 sky130_fd_sc_hd__xnor2_2 _32794_ (.A(_04515_),
    .B(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__a21oi_2 _32795_ (.A1(_04163_),
    .A2(_04168_),
    .B1(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__and3_2 _32796_ (.A(_04163_),
    .B(_04168_),
    .C(_04518_),
    .X(_04520_));
 sky130_fd_sc_hd__or2_2 _32797_ (.A(_04519_),
    .B(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__xor2_2 _32798_ (.A(_04513_),
    .B(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__a32oi_2 _32799_ (.A1(_04140_),
    .A2(_04146_),
    .A3(_04147_),
    .B1(_04149_),
    .B2(_04137_),
    .Y(_04523_));
 sky130_fd_sc_hd__xor2_2 _32800_ (.A(_04522_),
    .B(_04523_),
    .X(_04524_));
 sky130_fd_sc_hd__xor2_2 _32801_ (.A(_04512_),
    .B(_04524_),
    .X(_04525_));
 sky130_fd_sc_hd__o21a_2 _32802_ (.A1(_04492_),
    .A2(_04493_),
    .B1(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__nor3_2 _32803_ (.A(_04492_),
    .B(_04493_),
    .C(_04525_),
    .Y(_04528_));
 sky130_fd_sc_hd__nor2_2 _32804_ (.A(_04526_),
    .B(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__xnor2_2 _32805_ (.A(_04491_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__or2_2 _32806_ (.A(_04169_),
    .B(_04175_),
    .X(_04531_));
 sky130_fd_sc_hd__o21a_2 _32807_ (.A1(_04173_),
    .A2(_04174_),
    .B1(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__and4_2 _32808_ (.A(_01039_),
    .B(_14411_),
    .C(_00268_),
    .D(_01643_),
    .X(_04533_));
 sky130_fd_sc_hd__o22a_2 _32809_ (.A1(_01605_),
    .A2(_04162_),
    .B1(_01070_),
    .B2(_02608_),
    .X(_04534_));
 sky130_fd_sc_hd__nor2_2 _32810_ (.A(_04533_),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__nand2_2 _32811_ (.A(_03023_),
    .B(_04138_),
    .Y(_04536_));
 sky130_fd_sc_hd__xnor2_2 _32812_ (.A(_04535_),
    .B(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__and3_2 _32813_ (.A(_13544_),
    .B(_03438_),
    .C(_04170_),
    .X(_04539_));
 sky130_fd_sc_hd__and2_2 _32814_ (.A(_04171_),
    .B(_04172_),
    .X(_04540_));
 sky130_fd_sc_hd__and3_2 _32815_ (.A(_13544_),
    .B(_02641_),
    .C(_04170_),
    .X(_04541_));
 sky130_fd_sc_hd__o22a_2 _32816_ (.A1(_18791_),
    .A2(_01087_),
    .B1(_02389_),
    .B2(_14626_),
    .X(_04542_));
 sky130_fd_sc_hd__or2_2 _32817_ (.A(_04541_),
    .B(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__nand2_2 _32818_ (.A(_13889_),
    .B(_01650_),
    .Y(_04544_));
 sky130_fd_sc_hd__xor2_2 _32819_ (.A(_04543_),
    .B(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__o21ai_2 _32820_ (.A1(_04539_),
    .A2(_04540_),
    .B1(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__or3_2 _32821_ (.A(_04539_),
    .B(_04540_),
    .C(_04545_),
    .X(_04547_));
 sky130_fd_sc_hd__and2_2 _32822_ (.A(_04546_),
    .B(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__xor2_2 _32823_ (.A(_04537_),
    .B(_04548_),
    .X(_04550_));
 sky130_fd_sc_hd__xor2_2 _32824_ (.A(_04197_),
    .B(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__xor2_2 _32825_ (.A(_04532_),
    .B(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__and3_2 _32826_ (.A(_02626_),
    .B(_03994_),
    .C(_04195_),
    .X(_04553_));
 sky130_fd_sc_hd__a22o_2 _32827_ (.A1(_02626_),
    .A2(_03457_),
    .B1(_03454_),
    .B2(_14636_),
    .X(_04554_));
 sky130_fd_sc_hd__or3_2 _32828_ (.A(_12852_),
    .B(_02652_),
    .C(_04189_),
    .X(_04555_));
 sky130_fd_sc_hd__and2_2 _32829_ (.A(_04554_),
    .B(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__o21a_2 _32830_ (.A1(_04193_),
    .A2(_04553_),
    .B1(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__nor3_2 _32831_ (.A(_04193_),
    .B(_04553_),
    .C(_04556_),
    .Y(_04558_));
 sky130_fd_sc_hd__or2_2 _32832_ (.A(_04557_),
    .B(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__o2bb2a_2 _32833_ (.A1_N(_04182_),
    .A2_N(_04184_),
    .B1(_12823_),
    .B2(_03068_),
    .X(_04561_));
 sky130_fd_sc_hd__a2bb2o_2 _32834_ (.A1_N(_18368_),
    .A2_N(_04181_),
    .B1(_04005_),
    .B2(_18192_),
    .X(_04562_));
 sky130_fd_sc_hd__o21a_2 _32835_ (.A1(_13856_),
    .A2(_03068_),
    .B1(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__xnor2_2 _32836_ (.A(_04561_),
    .B(_04563_),
    .Y(_04564_));
 sky130_fd_sc_hd__xnor2_2 _32837_ (.A(_04559_),
    .B(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__nand2_2 _32838_ (.A(_04180_),
    .B(_04185_),
    .Y(_04566_));
 sky130_fd_sc_hd__nor2_2 _32839_ (.A(_04180_),
    .B(_04185_),
    .Y(_04567_));
 sky130_fd_sc_hd__a21oi_2 _32840_ (.A1(_04566_),
    .A2(_04200_),
    .B1(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__xnor2_2 _32841_ (.A(_04565_),
    .B(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__xnor2_2 _32842_ (.A(_04552_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__and2b_2 _32843_ (.A_N(_04203_),
    .B(_04201_),
    .X(_04572_));
 sky130_fd_sc_hd__a21oi_2 _32844_ (.A1(_04179_),
    .A2(_04204_),
    .B1(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__xnor2_2 _32845_ (.A(_04570_),
    .B(_04573_),
    .Y(_04574_));
 sky130_fd_sc_hd__xnor2_2 _32846_ (.A(_04530_),
    .B(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__and2b_2 _32847_ (.A_N(_04205_),
    .B(_04207_),
    .X(_04576_));
 sky130_fd_sc_hd__a21oi_2 _32848_ (.A1(_04157_),
    .A2(_04208_),
    .B1(_04576_),
    .Y(_04577_));
 sky130_fd_sc_hd__xor2_2 _32849_ (.A(_04575_),
    .B(_04577_),
    .X(_04578_));
 sky130_fd_sc_hd__xnor2_2 _32850_ (.A(_04489_),
    .B(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__nor2_2 _32851_ (.A(_04209_),
    .B(_04212_),
    .Y(_04580_));
 sky130_fd_sc_hd__a21oi_2 _32852_ (.A1(_04114_),
    .A2(_04213_),
    .B1(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__xor2_2 _32853_ (.A(_04579_),
    .B(_04581_),
    .X(_04583_));
 sky130_fd_sc_hd__xnor2_2 _32854_ (.A(_04441_),
    .B(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__nor2_2 _32855_ (.A(_04214_),
    .B(_04216_),
    .Y(_04585_));
 sky130_fd_sc_hd__a21oi_2 _32856_ (.A1(_04066_),
    .A2(_04217_),
    .B1(_04585_),
    .Y(_04586_));
 sky130_fd_sc_hd__xor2_2 _32857_ (.A(_04584_),
    .B(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__xnor2_2 _32858_ (.A(_04064_),
    .B(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__nor2_2 _32859_ (.A(_04218_),
    .B(_04220_),
    .Y(_04589_));
 sky130_fd_sc_hd__a21oi_2 _32860_ (.A1(_03879_),
    .A2(_04222_),
    .B1(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__xnor2_2 _32861_ (.A(_04588_),
    .B(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__a21o_2 _32862_ (.A1(_04226_),
    .A2(_04229_),
    .B1(_04591_),
    .X(_04592_));
 sky130_fd_sc_hd__nand3_2 _32863_ (.A(_04226_),
    .B(_04229_),
    .C(_04591_),
    .Y(_04594_));
 sky130_fd_sc_hd__and2b_2 _32864_ (.A_N(_04394_),
    .B(_04395_),
    .X(_04595_));
 sky130_fd_sc_hd__and2_2 _32865_ (.A(iY[39]),
    .B(iX[62]),
    .X(_04596_));
 sky130_fd_sc_hd__a21o_2 _32866_ (.A1(iY[38]),
    .A2(iX[63]),
    .B1(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__nand3_2 _32867_ (.A(iY[38]),
    .B(iX[63]),
    .C(_04596_),
    .Y(_04598_));
 sky130_fd_sc_hd__nand2_2 _32868_ (.A(_04597_),
    .B(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__nand2_2 _32869_ (.A(iY[40]),
    .B(iX[61]),
    .Y(_04600_));
 sky130_fd_sc_hd__xor2_2 _32870_ (.A(_04599_),
    .B(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__o21ai_2 _32871_ (.A1(_04240_),
    .A2(_04244_),
    .B1(_04601_),
    .Y(_04602_));
 sky130_fd_sc_hd__or3_2 _32872_ (.A(_04240_),
    .B(_04244_),
    .C(_04601_),
    .X(_04603_));
 sky130_fd_sc_hd__nand2_2 _32873_ (.A(_04602_),
    .B(_04603_),
    .Y(_04605_));
 sky130_fd_sc_hd__nand2_2 _32874_ (.A(_04250_),
    .B(_04605_),
    .Y(_04606_));
 sky130_fd_sc_hd__or2_2 _32875_ (.A(_04250_),
    .B(_04605_),
    .X(_04607_));
 sky130_fd_sc_hd__and2_2 _32876_ (.A(_04606_),
    .B(_04607_),
    .X(_04608_));
 sky130_fd_sc_hd__and2b_2 _32877_ (.A_N(_04271_),
    .B(_04270_),
    .X(_04609_));
 sky130_fd_sc_hd__or2b_2 _32878_ (.A(_04248_),
    .B_N(_04237_),
    .X(_04610_));
 sky130_fd_sc_hd__and4_2 _32879_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[56]),
    .D(iX[57]),
    .X(_04611_));
 sky130_fd_sc_hd__a22oi_2 _32880_ (.A1(iY[45]),
    .A2(iX[56]),
    .B1(iX[57]),
    .B2(iY[44]),
    .Y(_04612_));
 sky130_fd_sc_hd__nor2_2 _32881_ (.A(_04611_),
    .B(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__nand2_2 _32882_ (.A(iY[46]),
    .B(iX[55]),
    .Y(_04614_));
 sky130_fd_sc_hd__xnor2_2 _32883_ (.A(_04613_),
    .B(_04614_),
    .Y(_04616_));
 sky130_fd_sc_hd__and4_2 _32884_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[59]),
    .D(iX[60]),
    .X(_04617_));
 sky130_fd_sc_hd__a22oi_2 _32885_ (.A1(iY[42]),
    .A2(iX[59]),
    .B1(iX[60]),
    .B2(iY[41]),
    .Y(_04618_));
 sky130_fd_sc_hd__nor2_2 _32886_ (.A(_04617_),
    .B(_04618_),
    .Y(_04619_));
 sky130_fd_sc_hd__nand2_2 _32887_ (.A(iY[43]),
    .B(iX[58]),
    .Y(_04620_));
 sky130_fd_sc_hd__xnor2_2 _32888_ (.A(_04619_),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__o21ba_2 _32889_ (.A1(_04267_),
    .A2(_04269_),
    .B1_N(_04266_),
    .X(_04622_));
 sky130_fd_sc_hd__xnor2_2 _32890_ (.A(_04621_),
    .B(_04622_),
    .Y(_04623_));
 sky130_fd_sc_hd__and2_2 _32891_ (.A(_04616_),
    .B(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__nor2_2 _32892_ (.A(_04616_),
    .B(_04623_),
    .Y(_04625_));
 sky130_fd_sc_hd__or2_2 _32893_ (.A(_04624_),
    .B(_04625_),
    .X(_04627_));
 sky130_fd_sc_hd__a21o_2 _32894_ (.A1(_04246_),
    .A2(_04610_),
    .B1(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__nand3_2 _32895_ (.A(_04246_),
    .B(_04610_),
    .C(_04627_),
    .Y(_04629_));
 sky130_fd_sc_hd__o211ai_2 _32896_ (.A1(_04609_),
    .A2(_04273_),
    .B1(_04628_),
    .C1(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__a211o_2 _32897_ (.A1(_04628_),
    .A2(_04629_),
    .B1(_04609_),
    .C1(_04273_),
    .X(_04631_));
 sky130_fd_sc_hd__nand3_2 _32898_ (.A(_04608_),
    .B(_04630_),
    .C(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__a21oi_2 _32899_ (.A1(_04630_),
    .A2(_04631_),
    .B1(_04608_),
    .Y(_04633_));
 sky130_fd_sc_hd__inv_2 _32900_ (.A(_04633_),
    .Y(_04634_));
 sky130_fd_sc_hd__a31o_2 _32901_ (.A1(_04256_),
    .A2(_04279_),
    .A3(_04280_),
    .B1(_04255_),
    .X(_04635_));
 sky130_fd_sc_hd__and3_2 _32902_ (.A(_04632_),
    .B(_04634_),
    .C(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__a21oi_2 _32903_ (.A1(_04632_),
    .A2(_04634_),
    .B1(_04635_),
    .Y(_04638_));
 sky130_fd_sc_hd__nor2_2 _32904_ (.A(_04636_),
    .B(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__inv_2 _32905_ (.A(_04316_),
    .Y(_04640_));
 sky130_fd_sc_hd__and4_2 _32906_ (.A(iX[47]),
    .B(iX[48]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_04641_));
 sky130_fd_sc_hd__a22oi_2 _32907_ (.A1(iX[48]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[47]),
    .Y(_04642_));
 sky130_fd_sc_hd__nor2_2 _32908_ (.A(_04641_),
    .B(_04642_),
    .Y(_04643_));
 sky130_fd_sc_hd__nand2_2 _32909_ (.A(iX[46]),
    .B(iY[55]),
    .Y(_04644_));
 sky130_fd_sc_hd__xnor2_2 _32910_ (.A(_04643_),
    .B(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__and4_2 _32911_ (.A(iX[50]),
    .B(iY[50]),
    .C(iX[51]),
    .D(iY[51]),
    .X(_04646_));
 sky130_fd_sc_hd__a22oi_2 _32912_ (.A1(iY[50]),
    .A2(iX[51]),
    .B1(iY[51]),
    .B2(iX[50]),
    .Y(_04647_));
 sky130_fd_sc_hd__nor2_2 _32913_ (.A(_04646_),
    .B(_04647_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand2_2 _32914_ (.A(iX[49]),
    .B(iY[52]),
    .Y(_04650_));
 sky130_fd_sc_hd__xnor2_2 _32915_ (.A(_04649_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__o21ba_2 _32916_ (.A1(_04294_),
    .A2(_04296_),
    .B1_N(_04293_),
    .X(_04652_));
 sky130_fd_sc_hd__xnor2_2 _32917_ (.A(_04651_),
    .B(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__and2_2 _32918_ (.A(_04645_),
    .B(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__nor2_2 _32919_ (.A(_04645_),
    .B(_04653_),
    .Y(_04655_));
 sky130_fd_sc_hd__or2_2 _32920_ (.A(_04654_),
    .B(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__or3_2 _32921_ (.A(_04305_),
    .B(_04309_),
    .C(_04310_),
    .X(_04657_));
 sky130_fd_sc_hd__o21ba_2 _32922_ (.A1(_04261_),
    .A2(_04263_),
    .B1_N(_04260_),
    .X(_04658_));
 sky130_fd_sc_hd__and4_2 _32923_ (.A(iY[47]),
    .B(iY[48]),
    .C(iX[53]),
    .D(iX[54]),
    .X(_04660_));
 sky130_fd_sc_hd__a22oi_2 _32924_ (.A1(iY[48]),
    .A2(iX[53]),
    .B1(iX[54]),
    .B2(iY[47]),
    .Y(_04661_));
 sky130_fd_sc_hd__nand2_2 _32925_ (.A(iY[49]),
    .B(iX[52]),
    .Y(_04662_));
 sky130_fd_sc_hd__o21a_2 _32926_ (.A1(_04660_),
    .A2(_04661_),
    .B1(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__nor3_2 _32927_ (.A(_04660_),
    .B(_04661_),
    .C(_04662_),
    .Y(_04664_));
 sky130_fd_sc_hd__nor2_2 _32928_ (.A(_04663_),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__xnor2_2 _32929_ (.A(_04658_),
    .B(_04665_),
    .Y(_04666_));
 sky130_fd_sc_hd__o21ai_2 _32930_ (.A1(_04306_),
    .A2(_04310_),
    .B1(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__or3_2 _32931_ (.A(_04306_),
    .B(_04310_),
    .C(_04666_),
    .X(_04668_));
 sky130_fd_sc_hd__nand2_2 _32932_ (.A(_04667_),
    .B(_04668_),
    .Y(_04669_));
 sky130_fd_sc_hd__a21oi_2 _32933_ (.A1(_04657_),
    .A2(_04313_),
    .B1(_04669_),
    .Y(_04671_));
 sky130_fd_sc_hd__and3_2 _32934_ (.A(_04657_),
    .B(_04313_),
    .C(_04669_),
    .X(_04672_));
 sky130_fd_sc_hd__or3_2 _32935_ (.A(_04656_),
    .B(_04671_),
    .C(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__o21ai_2 _32936_ (.A1(_04671_),
    .A2(_04672_),
    .B1(_04656_),
    .Y(_04674_));
 sky130_fd_sc_hd__nand2_2 _32937_ (.A(_04673_),
    .B(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__a21oi_2 _32938_ (.A1(_04277_),
    .A2(_04279_),
    .B1(_04675_),
    .Y(_04676_));
 sky130_fd_sc_hd__and3_2 _32939_ (.A(_04277_),
    .B(_04279_),
    .C(_04675_),
    .X(_04677_));
 sky130_fd_sc_hd__a211oi_2 _32940_ (.A1(_04640_),
    .A2(_04318_),
    .B1(_04676_),
    .C1(_04677_),
    .Y(_04678_));
 sky130_fd_sc_hd__o211a_2 _32941_ (.A1(_04676_),
    .A2(_04677_),
    .B1(_04640_),
    .C1(_04318_),
    .X(_04679_));
 sky130_fd_sc_hd__nor2_2 _32942_ (.A(_04678_),
    .B(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__xnor2_2 _32943_ (.A(_04639_),
    .B(_04680_),
    .Y(_04682_));
 sky130_fd_sc_hd__o21ba_2 _32944_ (.A1(_04282_),
    .A2(_04283_),
    .B1_N(_04327_),
    .X(_04683_));
 sky130_fd_sc_hd__xnor2_2 _32945_ (.A(_04682_),
    .B(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__a21bo_2 _32946_ (.A1(_04351_),
    .A2(_04372_),
    .B1_N(_04371_),
    .X(_04685_));
 sky130_fd_sc_hd__and2_2 _32947_ (.A(_04285_),
    .B(_04324_),
    .X(_04686_));
 sky130_fd_sc_hd__or2b_2 _32948_ (.A(_04340_),
    .B_N(_04339_),
    .X(_04687_));
 sky130_fd_sc_hd__and4_2 _32949_ (.A(iX[41]),
    .B(iX[42]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_04688_));
 sky130_fd_sc_hd__a22oi_2 _32950_ (.A1(iX[42]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[41]),
    .Y(_04689_));
 sky130_fd_sc_hd__nor2_2 _32951_ (.A(_04688_),
    .B(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__nand2_2 _32952_ (.A(iX[40]),
    .B(iY[61]),
    .Y(_04691_));
 sky130_fd_sc_hd__xnor2_2 _32953_ (.A(_04690_),
    .B(_04691_),
    .Y(_04693_));
 sky130_fd_sc_hd__o21ba_2 _32954_ (.A1(_04336_),
    .A2(_04338_),
    .B1_N(_04335_),
    .X(_04694_));
 sky130_fd_sc_hd__xnor2_2 _32955_ (.A(_04693_),
    .B(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__and2_2 _32956_ (.A(iX[39]),
    .B(iY[62]),
    .X(_04696_));
 sky130_fd_sc_hd__or2_2 _32957_ (.A(_04695_),
    .B(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__nand2_2 _32958_ (.A(_04695_),
    .B(_04696_),
    .Y(_04698_));
 sky130_fd_sc_hd__nand2_2 _32959_ (.A(_04697_),
    .B(_04698_),
    .Y(_04699_));
 sky130_fd_sc_hd__a21oi_2 _32960_ (.A1(_04687_),
    .A2(_04345_),
    .B1(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__and3_2 _32961_ (.A(_04687_),
    .B(_04345_),
    .C(_04699_),
    .X(_04701_));
 sky130_fd_sc_hd__nor2_2 _32962_ (.A(_04700_),
    .B(_04701_),
    .Y(_04702_));
 sky130_fd_sc_hd__nand2_2 _32963_ (.A(iX[38]),
    .B(iY[63]),
    .Y(_04704_));
 sky130_fd_sc_hd__xnor2_2 _32964_ (.A(_04702_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__or2b_2 _32965_ (.A(_04357_),
    .B_N(_04362_),
    .X(_04706_));
 sky130_fd_sc_hd__or2b_2 _32966_ (.A(_04356_),
    .B_N(_04364_),
    .X(_04707_));
 sky130_fd_sc_hd__and2b_2 _32967_ (.A_N(_04299_),
    .B(_04297_),
    .X(_04708_));
 sky130_fd_sc_hd__o21ba_2 _32968_ (.A1(_04359_),
    .A2(_04361_),
    .B1_N(_04358_),
    .X(_04709_));
 sky130_fd_sc_hd__o21ba_2 _32969_ (.A1(_04289_),
    .A2(_04291_),
    .B1_N(_04288_),
    .X(_04710_));
 sky130_fd_sc_hd__and4_2 _32970_ (.A(iX[44]),
    .B(iX[45]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_04711_));
 sky130_fd_sc_hd__a22oi_2 _32971_ (.A1(iX[45]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[44]),
    .Y(_04712_));
 sky130_fd_sc_hd__nor2_2 _32972_ (.A(_04711_),
    .B(_04712_),
    .Y(_04713_));
 sky130_fd_sc_hd__nand2_2 _32973_ (.A(iX[43]),
    .B(iY[58]),
    .Y(_04715_));
 sky130_fd_sc_hd__xnor2_2 _32974_ (.A(_04713_),
    .B(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hd__xnor2_2 _32975_ (.A(_04710_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__xnor2_2 _32976_ (.A(_04709_),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__o21a_2 _32977_ (.A1(_04708_),
    .A2(_04301_),
    .B1(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__nor3_2 _32978_ (.A(_04708_),
    .B(_04301_),
    .C(_04718_),
    .Y(_04720_));
 sky130_fd_sc_hd__a211oi_2 _32979_ (.A1(_04706_),
    .A2(_04707_),
    .B1(_04719_),
    .C1(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__o211a_2 _32980_ (.A1(_04719_),
    .A2(_04720_),
    .B1(_04706_),
    .C1(_04707_),
    .X(_04722_));
 sky130_fd_sc_hd__nor2_2 _32981_ (.A(_04366_),
    .B(_04368_),
    .Y(_04723_));
 sky130_fd_sc_hd__or3_2 _32982_ (.A(_04721_),
    .B(_04722_),
    .C(_04723_),
    .X(_04724_));
 sky130_fd_sc_hd__o21ai_2 _32983_ (.A1(_04721_),
    .A2(_04722_),
    .B1(_04723_),
    .Y(_04726_));
 sky130_fd_sc_hd__and3_2 _32984_ (.A(_04705_),
    .B(_04724_),
    .C(_04726_),
    .X(_04727_));
 sky130_fd_sc_hd__a21oi_2 _32985_ (.A1(_04724_),
    .A2(_04726_),
    .B1(_04705_),
    .Y(_04728_));
 sky130_fd_sc_hd__nor2_2 _32986_ (.A(_04727_),
    .B(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hd__o21ai_2 _32987_ (.A1(_04322_),
    .A2(_04686_),
    .B1(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__or3_2 _32988_ (.A(_04322_),
    .B(_04686_),
    .C(_04729_),
    .X(_04731_));
 sky130_fd_sc_hd__and3_2 _32989_ (.A(_04685_),
    .B(_04730_),
    .C(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__a21oi_2 _32990_ (.A1(_04730_),
    .A2(_04731_),
    .B1(_04685_),
    .Y(_04733_));
 sky130_fd_sc_hd__nor2_2 _32991_ (.A(_04732_),
    .B(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__xor2_2 _32992_ (.A(_04684_),
    .B(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__a21o_2 _32993_ (.A1(_04329_),
    .A2(_04381_),
    .B1(_04735_),
    .X(_04737_));
 sky130_fd_sc_hd__nand3_2 _32994_ (.A(_04329_),
    .B(_04381_),
    .C(_04735_),
    .Y(_04738_));
 sky130_fd_sc_hd__and2_2 _32995_ (.A(_04737_),
    .B(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__o21ba_2 _32996_ (.A1(_04333_),
    .A2(_04378_),
    .B1_N(_04377_),
    .X(_04740_));
 sky130_fd_sc_hd__xnor2_2 _32997_ (.A(_04739_),
    .B(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__o21a_2 _32998_ (.A1(_04388_),
    .A2(_04390_),
    .B1(_04386_),
    .X(_04742_));
 sky130_fd_sc_hd__xnor2_2 _32999_ (.A(_04741_),
    .B(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__a31oi_2 _33000_ (.A1(iX[37]),
    .A2(iY[63]),
    .A3(_04348_),
    .B1(_04346_),
    .Y(_04744_));
 sky130_fd_sc_hd__xnor2_2 _33001_ (.A(_04743_),
    .B(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__nor3_2 _33002_ (.A(_04392_),
    .B(_04595_),
    .C(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__o21ai_2 _33003_ (.A1(_04392_),
    .A2(_04595_),
    .B1(_04745_),
    .Y(_04748_));
 sky130_fd_sc_hd__or2b_2 _33004_ (.A(_04746_),
    .B_N(_04748_),
    .X(_04749_));
 sky130_fd_sc_hd__a21bo_2 _33005_ (.A1(_04399_),
    .A2(_04405_),
    .B1_N(_04398_),
    .X(_04750_));
 sky130_fd_sc_hd__xor2_2 _33006_ (.A(_04749_),
    .B(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__a21o_2 _33007_ (.A1(_04592_),
    .A2(_04594_),
    .B1(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__nand3_2 _33008_ (.A(_04592_),
    .B(_04594_),
    .C(_04751_),
    .Y(_04753_));
 sky130_fd_sc_hd__nand3b_2 _33009_ (.A_N(_12448_),
    .B(_04752_),
    .C(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__a21bo_2 _33010_ (.A1(_04752_),
    .A2(_04753_),
    .B1_N(_12448_),
    .X(_04755_));
 sky130_fd_sc_hd__nand2_2 _33011_ (.A(_04754_),
    .B(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__a21oi_2 _33012_ (.A1(_04052_),
    .A2(_04410_),
    .B1(_04408_),
    .Y(_04757_));
 sky130_fd_sc_hd__nor2_2 _33013_ (.A(_04756_),
    .B(_04757_),
    .Y(_04759_));
 sky130_fd_sc_hd__and2_2 _33014_ (.A(_04756_),
    .B(_04757_),
    .X(_04760_));
 sky130_fd_sc_hd__or2_2 _33015_ (.A(_04759_),
    .B(_04760_),
    .X(_04761_));
 sky130_fd_sc_hd__o21ba_2 _33016_ (.A1(_04415_),
    .A2(_04422_),
    .B1_N(_04413_),
    .X(_04762_));
 sky130_fd_sc_hd__xnor2_2 _33017_ (.A(_04761_),
    .B(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__and2b_2 _33018_ (.A_N(_12521_),
    .B(_04763_),
    .X(_04764_));
 sky130_fd_sc_hd__and2b_2 _33019_ (.A_N(_04763_),
    .B(_12521_),
    .X(_04765_));
 sky130_fd_sc_hd__nor2_2 _33020_ (.A(_04764_),
    .B(_04765_),
    .Y(_04766_));
 sky130_fd_sc_hd__nor2_2 _33021_ (.A(_04424_),
    .B(_04432_),
    .Y(_04767_));
 sky130_fd_sc_hd__xnor2_2 _33022_ (.A(_04766_),
    .B(_04767_),
    .Y(oO[69]));
 sky130_fd_sc_hd__xnor2_2 _33023_ (.A(_13062_),
    .B(_12694_),
    .Y(_04769_));
 sky130_fd_sc_hd__or2b_2 _33024_ (.A(_04487_),
    .B_N(_04445_),
    .X(_04770_));
 sky130_fd_sc_hd__or2b_2 _33025_ (.A(_04488_),
    .B_N(_04443_),
    .X(_04771_));
 sky130_fd_sc_hd__and2b_2 _33026_ (.A_N(_04462_),
    .B(_04463_),
    .X(_04772_));
 sky130_fd_sc_hd__a21oi_2 _33027_ (.A1(_04446_),
    .A2(_04464_),
    .B1(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__a21oi_2 _33028_ (.A1(_04770_),
    .A2(_04771_),
    .B1(_04773_),
    .Y(_04774_));
 sky130_fd_sc_hd__and3_2 _33029_ (.A(_04770_),
    .B(_04771_),
    .C(_04773_),
    .X(_04775_));
 sky130_fd_sc_hd__nor2_2 _33030_ (.A(_04774_),
    .B(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__and2b_2 _33031_ (.A_N(_04485_),
    .B(_04481_),
    .X(_04777_));
 sky130_fd_sc_hd__a21o_2 _33032_ (.A1(_04465_),
    .A2(_04486_),
    .B1(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__a21o_2 _33033_ (.A1(_04491_),
    .A2(_04529_),
    .B1(_04526_),
    .X(_04780_));
 sky130_fd_sc_hd__buf_1 _33034_ (.A(_02928_),
    .X(_04781_));
 sky130_fd_sc_hd__inv_2 _33035_ (.A(_04781_),
    .Y(_04782_));
 sky130_fd_sc_hd__nor2_2 _33036_ (.A(_00990_),
    .B(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__a32o_2 _33037_ (.A1(_01564_),
    .A2(_04451_),
    .A3(_04449_),
    .B1(_04783_),
    .B2(_04447_),
    .X(_04784_));
 sky130_fd_sc_hd__or2_2 _33038_ (.A(_16288_),
    .B(_02316_),
    .X(_04785_));
 sky130_fd_sc_hd__a2bb2o_2 _33039_ (.A1_N(_00990_),
    .A2_N(_02317_),
    .B1(_01522_),
    .B2(_01785_),
    .X(_04786_));
 sky130_fd_sc_hd__o21ai_2 _33040_ (.A1(_04448_),
    .A2(_04785_),
    .B1(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__nand2_2 _33041_ (.A(_02338_),
    .B(_04451_),
    .Y(_04788_));
 sky130_fd_sc_hd__xor2_2 _33042_ (.A(_04787_),
    .B(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__or4_2 _33043_ (.A(_01576_),
    .B(_01583_),
    .C(_02940_),
    .D(_01512_),
    .X(_04791_));
 sky130_fd_sc_hd__a22o_2 _33044_ (.A1(_15888_),
    .A2(_01757_),
    .B1(_00566_),
    .B2(_18157_),
    .X(_04792_));
 sky130_fd_sc_hd__nand2_2 _33045_ (.A(_04791_),
    .B(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__nand2_2 _33046_ (.A(_00999_),
    .B(_01733_),
    .Y(_04794_));
 sky130_fd_sc_hd__xnor2_2 _33047_ (.A(_04793_),
    .B(_04794_),
    .Y(_04795_));
 sky130_fd_sc_hd__o21a_2 _33048_ (.A1(_04456_),
    .A2(_04457_),
    .B1(_04454_),
    .X(_04796_));
 sky130_fd_sc_hd__xor2_2 _33049_ (.A(_04795_),
    .B(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__nand2_2 _33050_ (.A(_04789_),
    .B(_04797_),
    .Y(_04798_));
 sky130_fd_sc_hd__or2_2 _33051_ (.A(_04789_),
    .B(_04797_),
    .X(_04799_));
 sky130_fd_sc_hd__nand2_2 _33052_ (.A(_04798_),
    .B(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__nor2_2 _33053_ (.A(_04458_),
    .B(_04459_),
    .Y(_04802_));
 sky130_fd_sc_hd__a21o_2 _33054_ (.A1(_04453_),
    .A2(_04460_),
    .B1(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__xnor2_2 _33055_ (.A(_04800_),
    .B(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__xnor2_2 _33056_ (.A(_04784_),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__and2_2 _33057_ (.A(_04471_),
    .B(_04478_),
    .X(_04806_));
 sky130_fd_sc_hd__a21oi_2 _33058_ (.A1(_04473_),
    .A2(_04477_),
    .B1(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__o21bai_2 _33059_ (.A1(_04499_),
    .A2(_04510_),
    .B1_N(_04509_),
    .Y(_04808_));
 sky130_fd_sc_hd__nor2_2 _33060_ (.A(_04097_),
    .B(_04474_),
    .Y(_04809_));
 sky130_fd_sc_hd__a31o_2 _33061_ (.A1(_15888_),
    .A2(_04469_),
    .A3(_04475_),
    .B1(_04809_),
    .X(_04810_));
 sky130_fd_sc_hd__nand2_2 _33062_ (.A(_04495_),
    .B(_04498_),
    .Y(_04811_));
 sky130_fd_sc_hd__nand2_2 _33063_ (.A(_02989_),
    .B(_18734_),
    .Y(_04813_));
 sky130_fd_sc_hd__or2_2 _33064_ (.A(_04474_),
    .B(_04813_),
    .X(_04814_));
 sky130_fd_sc_hd__a22o_2 _33065_ (.A1(_02989_),
    .A2(_18328_),
    .B1(_18734_),
    .B2(_02994_),
    .X(_04815_));
 sky130_fd_sc_hd__nand2_2 _33066_ (.A(_04814_),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__nand2_2 _33067_ (.A(_02983_),
    .B(_02956_),
    .Y(_04817_));
 sky130_fd_sc_hd__xnor2_2 _33068_ (.A(_04816_),
    .B(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__xnor2_2 _33069_ (.A(_04811_),
    .B(_04818_),
    .Y(_04819_));
 sky130_fd_sc_hd__xnor2_2 _33070_ (.A(_04810_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__xor2_2 _33071_ (.A(_04808_),
    .B(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__xnor2_2 _33072_ (.A(_04807_),
    .B(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__and2b_2 _33073_ (.A_N(_04479_),
    .B(_04468_),
    .X(_04824_));
 sky130_fd_sc_hd__and2b_2 _33074_ (.A_N(_04480_),
    .B(_04467_),
    .X(_04825_));
 sky130_fd_sc_hd__nor2_2 _33075_ (.A(_04824_),
    .B(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__xnor2_2 _33076_ (.A(_04822_),
    .B(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hd__xnor2_2 _33077_ (.A(_04805_),
    .B(_04827_),
    .Y(_04828_));
 sky130_fd_sc_hd__xor2_2 _33078_ (.A(_04780_),
    .B(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__xnor2_2 _33079_ (.A(_04778_),
    .B(_04829_),
    .Y(_04830_));
 sky130_fd_sc_hd__nor2_2 _33080_ (.A(_04522_),
    .B(_04523_),
    .Y(_04831_));
 sky130_fd_sc_hd__a21o_2 _33081_ (.A1(_04512_),
    .A2(_04524_),
    .B1(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__or2b_2 _33082_ (.A(_04197_),
    .B_N(_04550_),
    .X(_04833_));
 sky130_fd_sc_hd__or2_2 _33083_ (.A(_04532_),
    .B(_04551_),
    .X(_04835_));
 sky130_fd_sc_hd__or4_2 _33084_ (.A(_01828_),
    .B(_00255_),
    .C(_18363_),
    .D(_17409_),
    .X(_04836_));
 sky130_fd_sc_hd__buf_1 _33085_ (.A(_17006_),
    .X(_04837_));
 sky130_fd_sc_hd__a22o_2 _33086_ (.A1(_04837_),
    .A2(_17394_),
    .B1(_02984_),
    .B2(_01040_),
    .X(_04838_));
 sky130_fd_sc_hd__and2_2 _33087_ (.A(_04836_),
    .B(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__nor2_2 _33088_ (.A(_01832_),
    .B(_17628_),
    .Y(_04840_));
 sky130_fd_sc_hd__xnor2_2 _33089_ (.A(_04839_),
    .B(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__nor2_2 _33090_ (.A(_15835_),
    .B(_18200_),
    .Y(_04842_));
 sky130_fd_sc_hd__xor2_2 _33091_ (.A(_04500_),
    .B(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__nor2_2 _33092_ (.A(_16619_),
    .B(_00649_),
    .Y(_04844_));
 sky130_fd_sc_hd__xnor2_2 _33093_ (.A(_04843_),
    .B(_04844_),
    .Y(_04846_));
 sky130_fd_sc_hd__buf_1 _33094_ (.A(_16619_),
    .X(_04847_));
 sky130_fd_sc_hd__nand2_2 _33095_ (.A(_04125_),
    .B(_04500_),
    .Y(_04848_));
 sky130_fd_sc_hd__o31a_2 _33096_ (.A1(_04504_),
    .A2(_04847_),
    .A3(_04502_),
    .B1(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__nor2_2 _33097_ (.A(_04846_),
    .B(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__and2_2 _33098_ (.A(_04846_),
    .B(_04849_),
    .X(_04851_));
 sky130_fd_sc_hd__nor2_2 _33099_ (.A(_04850_),
    .B(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__xnor2_2 _33100_ (.A(_04841_),
    .B(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__and2b_2 _33101_ (.A_N(_04521_),
    .B(_04513_),
    .X(_04854_));
 sky130_fd_sc_hd__nand2_2 _33102_ (.A(_04141_),
    .B(_04514_),
    .Y(_04855_));
 sky130_fd_sc_hd__a21bo_2 _33103_ (.A1(_04515_),
    .A2(_04517_),
    .B1_N(_04855_),
    .X(_04857_));
 sky130_fd_sc_hd__a31o_2 _33104_ (.A1(_14606_),
    .A2(_01647_),
    .A3(_04535_),
    .B1(_04533_),
    .X(_04858_));
 sky130_fd_sc_hd__or4_2 _33105_ (.A(_15173_),
    .B(_15154_),
    .C(_01066_),
    .D(_00271_),
    .X(_04859_));
 sky130_fd_sc_hd__a22o_2 _33106_ (.A1(_15586_),
    .A2(_00662_),
    .B1(_01647_),
    .B2(_15617_),
    .X(_04860_));
 sky130_fd_sc_hd__nand2_2 _33107_ (.A(_04859_),
    .B(_04860_),
    .Y(_04861_));
 sky130_fd_sc_hd__buf_1 _33108_ (.A(_18443_),
    .X(_04862_));
 sky130_fd_sc_hd__nor2_2 _33109_ (.A(_03388_),
    .B(_04862_),
    .Y(_04863_));
 sky130_fd_sc_hd__xnor2_2 _33110_ (.A(_04861_),
    .B(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__xnor2_2 _33111_ (.A(_04858_),
    .B(_04864_),
    .Y(_04865_));
 sky130_fd_sc_hd__xnor2_2 _33112_ (.A(_04857_),
    .B(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hd__o21a_2 _33113_ (.A1(_04519_),
    .A2(_04854_),
    .B1(_04866_),
    .X(_04868_));
 sky130_fd_sc_hd__inv_2 _33114_ (.A(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__or3_2 _33115_ (.A(_04519_),
    .B(_04854_),
    .C(_04866_),
    .X(_04870_));
 sky130_fd_sc_hd__and3_2 _33116_ (.A(_04853_),
    .B(_04869_),
    .C(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__a21oi_2 _33117_ (.A1(_04869_),
    .A2(_04870_),
    .B1(_04853_),
    .Y(_04872_));
 sky130_fd_sc_hd__a211oi_2 _33118_ (.A1(_04833_),
    .A2(_04835_),
    .B1(_04871_),
    .C1(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__o211a_2 _33119_ (.A1(_04871_),
    .A2(_04872_),
    .B1(_04833_),
    .C1(_04835_),
    .X(_04874_));
 sky130_fd_sc_hd__nor2_2 _33120_ (.A(_04873_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__xor2_2 _33121_ (.A(_04832_),
    .B(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__nand2_2 _33122_ (.A(_04537_),
    .B(_04548_),
    .Y(_04877_));
 sky130_fd_sc_hd__nand2_2 _33123_ (.A(_14411_),
    .B(_02629_),
    .Y(_04879_));
 sky130_fd_sc_hd__or3_2 _33124_ (.A(_13972_),
    .B(_00674_),
    .C(_00675_),
    .X(_04880_));
 sky130_fd_sc_hd__xor2_2 _33125_ (.A(_04879_),
    .B(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__nor2_2 _33126_ (.A(_01028_),
    .B(_04162_),
    .Y(_04882_));
 sky130_fd_sc_hd__xnor2_2 _33127_ (.A(_04881_),
    .B(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__or4_2 _33128_ (.A(_14626_),
    .B(_18791_),
    .C(_02391_),
    .D(_02643_),
    .X(_04884_));
 sky130_fd_sc_hd__a22o_2 _33129_ (.A1(_13544_),
    .A2(_02641_),
    .B1(_03457_),
    .B2(_17463_),
    .X(_04885_));
 sky130_fd_sc_hd__nand2_2 _33130_ (.A(_04884_),
    .B(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__nor2_2 _33131_ (.A(_02613_),
    .B(_02647_),
    .Y(_04887_));
 sky130_fd_sc_hd__xnor2_2 _33132_ (.A(_04886_),
    .B(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__o21ba_2 _33133_ (.A1(_04543_),
    .A2(_04544_),
    .B1_N(_04541_),
    .X(_04890_));
 sky130_fd_sc_hd__xor2_2 _33134_ (.A(_04888_),
    .B(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__xor2_2 _33135_ (.A(_04883_),
    .B(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__xnor2_2 _33136_ (.A(_04557_),
    .B(_04892_),
    .Y(_04893_));
 sky130_fd_sc_hd__a21oi_2 _33137_ (.A1(_04546_),
    .A2(_04877_),
    .B1(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__and3_2 _33138_ (.A(_04546_),
    .B(_04877_),
    .C(_04893_),
    .X(_04895_));
 sky130_fd_sc_hd__nor2_2 _33139_ (.A(_04894_),
    .B(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__or2b_2 _33140_ (.A(_04559_),
    .B_N(_04564_),
    .X(_04897_));
 sky130_fd_sc_hd__inv_2 _33141_ (.A(_04562_),
    .Y(_04898_));
 sky130_fd_sc_hd__o22a_2 _33142_ (.A1(_13856_),
    .A2(_03068_),
    .B1(_04561_),
    .B2(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__buf_1 _33143_ (.A(_02663_),
    .X(_04901_));
 sky130_fd_sc_hd__o22a_2 _33144_ (.A1(_00195_),
    .A2(_04181_),
    .B1(_04901_),
    .B2(_12848_),
    .X(_04902_));
 sky130_fd_sc_hd__a21o_2 _33145_ (.A1(_14344_),
    .A2(_03064_),
    .B1(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__xor2_2 _33146_ (.A(_04899_),
    .B(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__buf_1 _33147_ (.A(_03454_),
    .X(_04905_));
 sky130_fd_sc_hd__and3_2 _33148_ (.A(_02626_),
    .B(_04905_),
    .C(_04189_),
    .X(_04906_));
 sky130_fd_sc_hd__xnor2_2 _33149_ (.A(_04904_),
    .B(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__xor2_2 _33150_ (.A(_04897_),
    .B(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__xnor2_2 _33151_ (.A(_04896_),
    .B(_04908_),
    .Y(_04909_));
 sky130_fd_sc_hd__and2b_2 _33152_ (.A_N(_04568_),
    .B(_04565_),
    .X(_04910_));
 sky130_fd_sc_hd__a21oi_2 _33153_ (.A1(_04552_),
    .A2(_04569_),
    .B1(_04910_),
    .Y(_04912_));
 sky130_fd_sc_hd__xor2_2 _33154_ (.A(_04909_),
    .B(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__xor2_2 _33155_ (.A(_04876_),
    .B(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__or2_2 _33156_ (.A(_04530_),
    .B(_04574_),
    .X(_04915_));
 sky130_fd_sc_hd__o21a_2 _33157_ (.A1(_04570_),
    .A2(_04573_),
    .B1(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__xnor2_2 _33158_ (.A(_04914_),
    .B(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hd__xnor2_2 _33159_ (.A(_04830_),
    .B(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__nor2_2 _33160_ (.A(_04575_),
    .B(_04577_),
    .Y(_04919_));
 sky130_fd_sc_hd__a21o_2 _33161_ (.A1(_04489_),
    .A2(_04578_),
    .B1(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__xnor2_2 _33162_ (.A(_04918_),
    .B(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__xnor2_2 _33163_ (.A(_04776_),
    .B(_04921_),
    .Y(_04923_));
 sky130_fd_sc_hd__nor2_2 _33164_ (.A(_04579_),
    .B(_04581_),
    .Y(_04924_));
 sky130_fd_sc_hd__a21oi_2 _33165_ (.A1(_04441_),
    .A2(_04583_),
    .B1(_04924_),
    .Y(_04925_));
 sky130_fd_sc_hd__xor2_2 _33166_ (.A(_04923_),
    .B(_04925_),
    .X(_04926_));
 sky130_fd_sc_hd__xnor2_2 _33167_ (.A(_04438_),
    .B(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__nor2_2 _33168_ (.A(_04584_),
    .B(_04586_),
    .Y(_04928_));
 sky130_fd_sc_hd__a21oi_2 _33169_ (.A1(_04064_),
    .A2(_04587_),
    .B1(_04928_),
    .Y(_04929_));
 sky130_fd_sc_hd__xnor2_2 _33170_ (.A(_04927_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__or2_2 _33171_ (.A(_04228_),
    .B(_04591_),
    .X(_04931_));
 sky130_fd_sc_hd__a21o_2 _33172_ (.A1(_04055_),
    .A2(_04059_),
    .B1(_04931_),
    .X(_04932_));
 sky130_fd_sc_hd__a211o_2 _33173_ (.A1(_04588_),
    .A2(_04590_),
    .B1(_04223_),
    .C1(_04225_),
    .X(_04934_));
 sky130_fd_sc_hd__o21a_2 _33174_ (.A1(_04588_),
    .A2(_04590_),
    .B1(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__nand2_2 _33175_ (.A(_04932_),
    .B(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__xor2_2 _33176_ (.A(_04930_),
    .B(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__or2b_2 _33177_ (.A(_04740_),
    .B_N(_04739_),
    .X(_04938_));
 sky130_fd_sc_hd__inv_2 _33178_ (.A(_04671_),
    .Y(_04939_));
 sky130_fd_sc_hd__and4_2 _33179_ (.A(iX[48]),
    .B(iX[49]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_04940_));
 sky130_fd_sc_hd__a22oi_2 _33180_ (.A1(iX[49]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[48]),
    .Y(_04941_));
 sky130_fd_sc_hd__nor2_2 _33181_ (.A(_04940_),
    .B(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hd__nand2_2 _33182_ (.A(iX[47]),
    .B(iY[55]),
    .Y(_04943_));
 sky130_fd_sc_hd__xnor2_2 _33183_ (.A(_04942_),
    .B(_04943_),
    .Y(_04945_));
 sky130_fd_sc_hd__and4_2 _33184_ (.A(iY[50]),
    .B(iX[51]),
    .C(iY[51]),
    .D(iX[52]),
    .X(_04946_));
 sky130_fd_sc_hd__a22oi_2 _33185_ (.A1(iX[51]),
    .A2(iY[51]),
    .B1(iX[52]),
    .B2(iY[50]),
    .Y(_04947_));
 sky130_fd_sc_hd__nor2_2 _33186_ (.A(_04946_),
    .B(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__nand2_2 _33187_ (.A(iX[50]),
    .B(iY[52]),
    .Y(_04949_));
 sky130_fd_sc_hd__xnor2_2 _33188_ (.A(_04948_),
    .B(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__o21ba_2 _33189_ (.A1(_04647_),
    .A2(_04650_),
    .B1_N(_04646_),
    .X(_04951_));
 sky130_fd_sc_hd__xnor2_2 _33190_ (.A(_04950_),
    .B(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__and2_2 _33191_ (.A(_04945_),
    .B(_04952_),
    .X(_04953_));
 sky130_fd_sc_hd__nor2_2 _33192_ (.A(_04945_),
    .B(_04952_),
    .Y(_04954_));
 sky130_fd_sc_hd__or2_2 _33193_ (.A(_04953_),
    .B(_04954_),
    .X(_04956_));
 sky130_fd_sc_hd__or3_2 _33194_ (.A(_04658_),
    .B(_04663_),
    .C(_04664_),
    .X(_04957_));
 sky130_fd_sc_hd__o21ba_2 _33195_ (.A1(_04612_),
    .A2(_04614_),
    .B1_N(_04611_),
    .X(_04958_));
 sky130_fd_sc_hd__and4_2 _33196_ (.A(iY[47]),
    .B(iY[48]),
    .C(iX[54]),
    .D(iX[55]),
    .X(_04959_));
 sky130_fd_sc_hd__a22oi_2 _33197_ (.A1(iY[48]),
    .A2(iX[54]),
    .B1(iX[55]),
    .B2(iY[47]),
    .Y(_04960_));
 sky130_fd_sc_hd__nand2_2 _33198_ (.A(iY[49]),
    .B(iX[53]),
    .Y(_04961_));
 sky130_fd_sc_hd__o21a_2 _33199_ (.A1(_04959_),
    .A2(_04960_),
    .B1(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__nor3_2 _33200_ (.A(_04959_),
    .B(_04960_),
    .C(_04961_),
    .Y(_04963_));
 sky130_fd_sc_hd__nor2_2 _33201_ (.A(_04962_),
    .B(_04963_),
    .Y(_04964_));
 sky130_fd_sc_hd__xnor2_2 _33202_ (.A(_04958_),
    .B(_04964_),
    .Y(_04965_));
 sky130_fd_sc_hd__o21ai_2 _33203_ (.A1(_04660_),
    .A2(_04664_),
    .B1(_04965_),
    .Y(_04967_));
 sky130_fd_sc_hd__or3_2 _33204_ (.A(_04660_),
    .B(_04664_),
    .C(_04965_),
    .X(_04968_));
 sky130_fd_sc_hd__nand2_2 _33205_ (.A(_04967_),
    .B(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__a21oi_2 _33206_ (.A1(_04957_),
    .A2(_04667_),
    .B1(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__and3_2 _33207_ (.A(_04957_),
    .B(_04667_),
    .C(_04969_),
    .X(_04971_));
 sky130_fd_sc_hd__or3_2 _33208_ (.A(_04956_),
    .B(_04970_),
    .C(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__o21ai_2 _33209_ (.A1(_04970_),
    .A2(_04971_),
    .B1(_04956_),
    .Y(_04973_));
 sky130_fd_sc_hd__nand2_2 _33210_ (.A(_04972_),
    .B(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__a21oi_2 _33211_ (.A1(_04628_),
    .A2(_04630_),
    .B1(_04974_),
    .Y(_04975_));
 sky130_fd_sc_hd__and3_2 _33212_ (.A(_04628_),
    .B(_04630_),
    .C(_04974_),
    .X(_04976_));
 sky130_fd_sc_hd__a211oi_2 _33213_ (.A1(_04939_),
    .A2(_04673_),
    .B1(_04975_),
    .C1(_04976_),
    .Y(_04978_));
 sky130_fd_sc_hd__o211a_2 _33214_ (.A1(_04975_),
    .A2(_04976_),
    .B1(_04939_),
    .C1(_04673_),
    .X(_04979_));
 sky130_fd_sc_hd__nand2_2 _33215_ (.A(iY[40]),
    .B(iX[63]),
    .Y(_04980_));
 sky130_fd_sc_hd__a22o_2 _33216_ (.A1(iY[40]),
    .A2(iX[62]),
    .B1(iX[63]),
    .B2(iY[39]),
    .X(_04981_));
 sky130_fd_sc_hd__o21a_2 _33217_ (.A1(_04239_),
    .A2(_04980_),
    .B1(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__o21ai_2 _33218_ (.A1(_04599_),
    .A2(_04600_),
    .B1(_04598_),
    .Y(_04983_));
 sky130_fd_sc_hd__nand2_2 _33219_ (.A(_04982_),
    .B(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__or2_2 _33220_ (.A(_04982_),
    .B(_04983_),
    .X(_04985_));
 sky130_fd_sc_hd__and2_2 _33221_ (.A(_04984_),
    .B(_04985_),
    .X(_04986_));
 sky130_fd_sc_hd__and2b_2 _33222_ (.A_N(_04622_),
    .B(_04621_),
    .X(_04987_));
 sky130_fd_sc_hd__and4_2 _33223_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[57]),
    .D(iX[58]),
    .X(_04989_));
 sky130_fd_sc_hd__a22oi_2 _33224_ (.A1(iY[45]),
    .A2(iX[57]),
    .B1(iX[58]),
    .B2(iY[44]),
    .Y(_04990_));
 sky130_fd_sc_hd__nor2_2 _33225_ (.A(_04989_),
    .B(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__nand2_2 _33226_ (.A(iY[46]),
    .B(iX[56]),
    .Y(_04992_));
 sky130_fd_sc_hd__xnor2_2 _33227_ (.A(_04991_),
    .B(_04992_),
    .Y(_04993_));
 sky130_fd_sc_hd__and4_2 _33228_ (.A(iY[41]),
    .B(iY[42]),
    .C(iX[60]),
    .D(iX[61]),
    .X(_04994_));
 sky130_fd_sc_hd__a22oi_2 _33229_ (.A1(iY[42]),
    .A2(iX[60]),
    .B1(iX[61]),
    .B2(iY[41]),
    .Y(_04995_));
 sky130_fd_sc_hd__nor2_2 _33230_ (.A(_04994_),
    .B(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand2_2 _33231_ (.A(iY[43]),
    .B(iX[59]),
    .Y(_04997_));
 sky130_fd_sc_hd__xnor2_2 _33232_ (.A(_04996_),
    .B(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__o21ba_2 _33233_ (.A1(_04618_),
    .A2(_04620_),
    .B1_N(_04617_),
    .X(_05000_));
 sky130_fd_sc_hd__xnor2_2 _33234_ (.A(_04998_),
    .B(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__xnor2_2 _33235_ (.A(_04993_),
    .B(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__or2_2 _33236_ (.A(_04602_),
    .B(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__nand2_2 _33237_ (.A(_04602_),
    .B(_05002_),
    .Y(_05004_));
 sky130_fd_sc_hd__and2_2 _33238_ (.A(_05003_),
    .B(_05004_),
    .X(_05005_));
 sky130_fd_sc_hd__o21ai_2 _33239_ (.A1(_04987_),
    .A2(_04624_),
    .B1(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__or3_2 _33240_ (.A(_04987_),
    .B(_04624_),
    .C(_05005_),
    .X(_05007_));
 sky130_fd_sc_hd__and3_2 _33241_ (.A(_04986_),
    .B(_05006_),
    .C(_05007_),
    .X(_05008_));
 sky130_fd_sc_hd__a21oi_2 _33242_ (.A1(_05006_),
    .A2(_05007_),
    .B1(_04986_),
    .Y(_05009_));
 sky130_fd_sc_hd__a211o_2 _33243_ (.A1(_04607_),
    .A2(_04632_),
    .B1(_05008_),
    .C1(_05009_),
    .X(_05011_));
 sky130_fd_sc_hd__o211ai_2 _33244_ (.A1(_05008_),
    .A2(_05009_),
    .B1(_04607_),
    .C1(_04632_),
    .Y(_05012_));
 sky130_fd_sc_hd__nand2_2 _33245_ (.A(_05011_),
    .B(_05012_),
    .Y(_05013_));
 sky130_fd_sc_hd__o21a_2 _33246_ (.A1(_04978_),
    .A2(_04979_),
    .B1(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__or3_2 _33247_ (.A(_05013_),
    .B(_04978_),
    .C(_04979_),
    .X(_05015_));
 sky130_fd_sc_hd__and2b_2 _33248_ (.A_N(_05014_),
    .B(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__a21o_2 _33249_ (.A1(_04639_),
    .A2(_04680_),
    .B1(_04636_),
    .X(_05017_));
 sky130_fd_sc_hd__xnor2_2 _33250_ (.A(_05016_),
    .B(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__a21boi_2 _33251_ (.A1(_04705_),
    .A2(_04726_),
    .B1_N(_04724_),
    .Y(_05019_));
 sky130_fd_sc_hd__or2b_2 _33252_ (.A(_04694_),
    .B_N(_04693_),
    .X(_05020_));
 sky130_fd_sc_hd__and4_2 _33253_ (.A(iX[42]),
    .B(iX[43]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_05022_));
 sky130_fd_sc_hd__a22oi_2 _33254_ (.A1(iX[43]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[42]),
    .Y(_05023_));
 sky130_fd_sc_hd__nor2_2 _33255_ (.A(_05022_),
    .B(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__nand2_2 _33256_ (.A(iX[41]),
    .B(iY[61]),
    .Y(_05025_));
 sky130_fd_sc_hd__xnor2_2 _33257_ (.A(_05024_),
    .B(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__o21ba_2 _33258_ (.A1(_04689_),
    .A2(_04691_),
    .B1_N(_04688_),
    .X(_05027_));
 sky130_fd_sc_hd__xnor2_2 _33259_ (.A(_05026_),
    .B(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__and2_2 _33260_ (.A(iX[40]),
    .B(iY[62]),
    .X(_05029_));
 sky130_fd_sc_hd__or2_2 _33261_ (.A(_05028_),
    .B(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__nand2_2 _33262_ (.A(_05028_),
    .B(_05029_),
    .Y(_05031_));
 sky130_fd_sc_hd__nand2_2 _33263_ (.A(_05030_),
    .B(_05031_),
    .Y(_05033_));
 sky130_fd_sc_hd__a21oi_2 _33264_ (.A1(_05020_),
    .A2(_04698_),
    .B1(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hd__and3_2 _33265_ (.A(_05020_),
    .B(_04698_),
    .C(_05033_),
    .X(_05035_));
 sky130_fd_sc_hd__nor2_2 _33266_ (.A(_05034_),
    .B(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__nand2_2 _33267_ (.A(iX[39]),
    .B(iY[63]),
    .Y(_05037_));
 sky130_fd_sc_hd__xnor2_2 _33268_ (.A(_05036_),
    .B(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__or2b_2 _33269_ (.A(_04710_),
    .B_N(_04716_),
    .X(_05039_));
 sky130_fd_sc_hd__or2b_2 _33270_ (.A(_04709_),
    .B_N(_04717_),
    .X(_05040_));
 sky130_fd_sc_hd__and2b_2 _33271_ (.A_N(_04652_),
    .B(_04651_),
    .X(_05041_));
 sky130_fd_sc_hd__o21ba_2 _33272_ (.A1(_04712_),
    .A2(_04715_),
    .B1_N(_04711_),
    .X(_05042_));
 sky130_fd_sc_hd__o21ba_2 _33273_ (.A1(_04642_),
    .A2(_04644_),
    .B1_N(_04641_),
    .X(_05044_));
 sky130_fd_sc_hd__and4_2 _33274_ (.A(iX[45]),
    .B(iX[46]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_05045_));
 sky130_fd_sc_hd__a22oi_2 _33275_ (.A1(iX[46]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[45]),
    .Y(_05046_));
 sky130_fd_sc_hd__nor2_2 _33276_ (.A(_05045_),
    .B(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__nand2_2 _33277_ (.A(iX[44]),
    .B(iY[58]),
    .Y(_05048_));
 sky130_fd_sc_hd__xnor2_2 _33278_ (.A(_05047_),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__xnor2_2 _33279_ (.A(_05044_),
    .B(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__xnor2_2 _33280_ (.A(_05042_),
    .B(_05050_),
    .Y(_05051_));
 sky130_fd_sc_hd__o21a_2 _33281_ (.A1(_05041_),
    .A2(_04654_),
    .B1(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__nor3_2 _33282_ (.A(_05041_),
    .B(_04654_),
    .C(_05051_),
    .Y(_05053_));
 sky130_fd_sc_hd__a211oi_2 _33283_ (.A1(_05039_),
    .A2(_05040_),
    .B1(_05052_),
    .C1(_05053_),
    .Y(_05055_));
 sky130_fd_sc_hd__o211a_2 _33284_ (.A1(_05052_),
    .A2(_05053_),
    .B1(_05039_),
    .C1(_05040_),
    .X(_05056_));
 sky130_fd_sc_hd__nor2_2 _33285_ (.A(_04719_),
    .B(_04721_),
    .Y(_05057_));
 sky130_fd_sc_hd__or3_2 _33286_ (.A(_05055_),
    .B(_05056_),
    .C(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__o21ai_2 _33287_ (.A1(_05055_),
    .A2(_05056_),
    .B1(_05057_),
    .Y(_05059_));
 sky130_fd_sc_hd__and3_2 _33288_ (.A(_05038_),
    .B(_05058_),
    .C(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__a21oi_2 _33289_ (.A1(_05058_),
    .A2(_05059_),
    .B1(_05038_),
    .Y(_05061_));
 sky130_fd_sc_hd__nor2_2 _33290_ (.A(_05060_),
    .B(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__o21ai_2 _33291_ (.A1(_04676_),
    .A2(_04678_),
    .B1(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__or3_2 _33292_ (.A(_04676_),
    .B(_04678_),
    .C(_05062_),
    .X(_05064_));
 sky130_fd_sc_hd__nand2_2 _33293_ (.A(_05063_),
    .B(_05064_),
    .Y(_05066_));
 sky130_fd_sc_hd__xnor2_2 _33294_ (.A(_05019_),
    .B(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__or2_2 _33295_ (.A(_05018_),
    .B(_05067_),
    .X(_05068_));
 sky130_fd_sc_hd__nand2_2 _33296_ (.A(_05018_),
    .B(_05067_),
    .Y(_05069_));
 sky130_fd_sc_hd__nand2_2 _33297_ (.A(_05068_),
    .B(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__and2b_2 _33298_ (.A_N(_04684_),
    .B(_04734_),
    .X(_05071_));
 sky130_fd_sc_hd__o21ba_2 _33299_ (.A1(_04682_),
    .A2(_04683_),
    .B1_N(_05071_),
    .X(_05072_));
 sky130_fd_sc_hd__xnor2_2 _33300_ (.A(_05070_),
    .B(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__a21bo_2 _33301_ (.A1(_04685_),
    .A2(_04731_),
    .B1_N(_04730_),
    .X(_05074_));
 sky130_fd_sc_hd__xor2_2 _33302_ (.A(_05073_),
    .B(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__a21o_2 _33303_ (.A1(_04737_),
    .A2(_04938_),
    .B1(_05075_),
    .X(_05077_));
 sky130_fd_sc_hd__nand3_2 _33304_ (.A(_04737_),
    .B(_04938_),
    .C(_05075_),
    .Y(_05078_));
 sky130_fd_sc_hd__nand2_2 _33305_ (.A(_05077_),
    .B(_05078_),
    .Y(_05079_));
 sky130_fd_sc_hd__a31o_2 _33306_ (.A1(iX[38]),
    .A2(iY[63]),
    .A3(_04702_),
    .B1(_04700_),
    .X(_05080_));
 sky130_fd_sc_hd__xor2_2 _33307_ (.A(_05079_),
    .B(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__or2b_2 _33308_ (.A(_04742_),
    .B_N(_04741_),
    .X(_05082_));
 sky130_fd_sc_hd__or2b_2 _33309_ (.A(_04744_),
    .B_N(_04743_),
    .X(_05083_));
 sky130_fd_sc_hd__nand2_2 _33310_ (.A(_05082_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__xor2_2 _33311_ (.A(_05081_),
    .B(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__a211o_2 _33312_ (.A1(_04402_),
    .A2(_04404_),
    .B1(_04749_),
    .C1(_04400_),
    .X(_05086_));
 sky130_fd_sc_hd__o21a_2 _33313_ (.A1(_04398_),
    .A2(_04746_),
    .B1(_04748_),
    .X(_05088_));
 sky130_fd_sc_hd__and2_2 _33314_ (.A(_05086_),
    .B(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__xor2_2 _33315_ (.A(_05085_),
    .B(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__inv_2 _33316_ (.A(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__xnor2_2 _33317_ (.A(_04937_),
    .B(_05091_),
    .Y(_05092_));
 sky130_fd_sc_hd__xnor2_2 _33318_ (.A(_04769_),
    .B(_05092_),
    .Y(_05093_));
 sky130_fd_sc_hd__and2_2 _33319_ (.A(_04753_),
    .B(_04754_),
    .X(_05094_));
 sky130_fd_sc_hd__xor2_2 _33320_ (.A(_05093_),
    .B(_05094_),
    .X(_05095_));
 sky130_fd_sc_hd__o21bai_2 _33321_ (.A1(_04413_),
    .A2(_04759_),
    .B1_N(_04760_),
    .Y(_05096_));
 sky130_fd_sc_hd__o31ai_2 _33322_ (.A1(_04415_),
    .A2(_04422_),
    .A3(_04761_),
    .B1(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__xor2_2 _33323_ (.A(_05095_),
    .B(_05097_),
    .X(_05099_));
 sky130_fd_sc_hd__nand2_2 _33324_ (.A(_12738_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__or2_2 _33325_ (.A(_12738_),
    .B(_05099_),
    .X(_05101_));
 sky130_fd_sc_hd__nand2_2 _33326_ (.A(_05100_),
    .B(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__or2b_2 _33327_ (.A(_12521_),
    .B_N(_04763_),
    .X(_05103_));
 sky130_fd_sc_hd__a21o_2 _33328_ (.A1(_04424_),
    .A2(_05103_),
    .B1(_04765_),
    .X(_05104_));
 sky130_fd_sc_hd__a21oi_2 _33329_ (.A1(_04432_),
    .A2(_04766_),
    .B1(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__xor2_2 _33330_ (.A(_05102_),
    .B(_05105_),
    .X(oO[70]));
 sky130_fd_sc_hd__nor2_2 _33331_ (.A(_05093_),
    .B(_05094_),
    .Y(_05106_));
 sky130_fd_sc_hd__a21oi_2 _33332_ (.A1(_05095_),
    .A2(_05097_),
    .B1(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__or2_2 _33333_ (.A(_04927_),
    .B(_04929_),
    .X(_05109_));
 sky130_fd_sc_hd__a21o_2 _33334_ (.A1(_04932_),
    .A2(_04935_),
    .B1(_04930_),
    .X(_05110_));
 sky130_fd_sc_hd__nor2_2 _33335_ (.A(_04923_),
    .B(_04925_),
    .Y(_05111_));
 sky130_fd_sc_hd__a21oi_2 _33336_ (.A1(_04438_),
    .A2(_04926_),
    .B1(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__or2b_2 _33337_ (.A(_04828_),
    .B_N(_04780_),
    .X(_05113_));
 sky130_fd_sc_hd__or2b_2 _33338_ (.A(_04829_),
    .B_N(_04778_),
    .X(_05114_));
 sky130_fd_sc_hd__a32oi_2 _33339_ (.A1(_04798_),
    .A2(_04799_),
    .A3(_04803_),
    .B1(_04804_),
    .B2(_04784_),
    .Y(_05115_));
 sky130_fd_sc_hd__a21oi_2 _33340_ (.A1(_05113_),
    .A2(_05114_),
    .B1(_05115_),
    .Y(_05116_));
 sky130_fd_sc_hd__and3_2 _33341_ (.A(_05113_),
    .B(_05114_),
    .C(_05115_),
    .X(_05117_));
 sky130_fd_sc_hd__nor2_2 _33342_ (.A(_05116_),
    .B(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__or2_2 _33343_ (.A(_04805_),
    .B(_04827_),
    .X(_05120_));
 sky130_fd_sc_hd__o21a_2 _33344_ (.A1(_04822_),
    .A2(_04826_),
    .B1(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__a21oi_2 _33345_ (.A1(_04832_),
    .A2(_04875_),
    .B1(_04873_),
    .Y(_05122_));
 sky130_fd_sc_hd__o22ai_2 _33346_ (.A1(_04448_),
    .A2(_04785_),
    .B1(_04787_),
    .B2(_04788_),
    .Y(_05123_));
 sky130_fd_sc_hd__nand2_2 _33347_ (.A(_00999_),
    .B(_01522_),
    .Y(_05124_));
 sky130_fd_sc_hd__xnor2_2 _33348_ (.A(_04785_),
    .B(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__nor2_2 _33349_ (.A(_00990_),
    .B(_03318_),
    .Y(_05126_));
 sky130_fd_sc_hd__xnor2_2 _33350_ (.A(_05125_),
    .B(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__or4_2 _33351_ (.A(_01583_),
    .B(_02463_),
    .C(_02940_),
    .D(_01512_),
    .X(_05128_));
 sky130_fd_sc_hd__a22o_2 _33352_ (.A1(_02983_),
    .A2(_01757_),
    .B1(_00566_),
    .B2(_15888_),
    .X(_05129_));
 sky130_fd_sc_hd__nand2_2 _33353_ (.A(_05128_),
    .B(_05129_),
    .Y(_05131_));
 sky130_fd_sc_hd__nand2_2 _33354_ (.A(_18157_),
    .B(_01733_),
    .Y(_05132_));
 sky130_fd_sc_hd__xnor2_2 _33355_ (.A(_05131_),
    .B(_05132_),
    .Y(_05133_));
 sky130_fd_sc_hd__o21a_2 _33356_ (.A1(_04793_),
    .A2(_04794_),
    .B1(_04791_),
    .X(_05134_));
 sky130_fd_sc_hd__xor2_2 _33357_ (.A(_05133_),
    .B(_05134_),
    .X(_05135_));
 sky130_fd_sc_hd__nand2_2 _33358_ (.A(_05127_),
    .B(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__or2_2 _33359_ (.A(_05127_),
    .B(_05135_),
    .X(_05137_));
 sky130_fd_sc_hd__nand2_2 _33360_ (.A(_05136_),
    .B(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__o21ai_2 _33361_ (.A1(_04795_),
    .A2(_04796_),
    .B1(_04798_),
    .Y(_05139_));
 sky130_fd_sc_hd__xnor2_2 _33362_ (.A(_05138_),
    .B(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__xnor2_2 _33363_ (.A(_05123_),
    .B(_05140_),
    .Y(_05142_));
 sky130_fd_sc_hd__or2b_2 _33364_ (.A(_04818_),
    .B_N(_04811_),
    .X(_05143_));
 sky130_fd_sc_hd__nand2_2 _33365_ (.A(_04810_),
    .B(_04819_),
    .Y(_05144_));
 sky130_fd_sc_hd__or2_2 _33366_ (.A(_04846_),
    .B(_04849_),
    .X(_05145_));
 sky130_fd_sc_hd__o21ai_2 _33367_ (.A1(_04841_),
    .A2(_04851_),
    .B1(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__o21ai_2 _33368_ (.A1(_04816_),
    .A2(_04817_),
    .B1(_04814_),
    .Y(_05147_));
 sky130_fd_sc_hd__a21bo_2 _33369_ (.A1(_04838_),
    .A2(_04840_),
    .B1_N(_04836_),
    .X(_05148_));
 sky130_fd_sc_hd__or3_2 _33370_ (.A(_01832_),
    .B(_18111_),
    .C(_18113_),
    .X(_05149_));
 sky130_fd_sc_hd__xor2_2 _33371_ (.A(_04813_),
    .B(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__nand2_2 _33372_ (.A(_02994_),
    .B(_02956_),
    .Y(_05151_));
 sky130_fd_sc_hd__xor2_2 _33373_ (.A(_05150_),
    .B(_05151_),
    .X(_05153_));
 sky130_fd_sc_hd__xor2_2 _33374_ (.A(_05148_),
    .B(_05153_),
    .X(_05154_));
 sky130_fd_sc_hd__xnor2_2 _33375_ (.A(_05147_),
    .B(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__xnor2_2 _33376_ (.A(_05146_),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__a21oi_2 _33377_ (.A1(_05143_),
    .A2(_05144_),
    .B1(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__and3_2 _33378_ (.A(_05143_),
    .B(_05144_),
    .C(_05156_),
    .X(_05158_));
 sky130_fd_sc_hd__nor2_2 _33379_ (.A(_05157_),
    .B(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__or2b_2 _33380_ (.A(_04820_),
    .B_N(_04808_),
    .X(_05160_));
 sky130_fd_sc_hd__o21a_2 _33381_ (.A1(_04807_),
    .A2(_04821_),
    .B1(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__xnor2_2 _33382_ (.A(_05159_),
    .B(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__xnor2_2 _33383_ (.A(_05142_),
    .B(_05162_),
    .Y(_05164_));
 sky130_fd_sc_hd__xnor2_2 _33384_ (.A(_05122_),
    .B(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__xnor2_2 _33385_ (.A(_05121_),
    .B(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__a21oi_2 _33386_ (.A1(_04557_),
    .A2(_04892_),
    .B1(_04894_),
    .Y(_05167_));
 sky130_fd_sc_hd__or4_2 _33387_ (.A(_00255_),
    .B(_00649_),
    .C(_18363_),
    .D(_17409_),
    .X(_05168_));
 sky130_fd_sc_hd__a22o_2 _33388_ (.A1(_01837_),
    .A2(_17394_),
    .B1(_02984_),
    .B2(_04837_),
    .X(_05169_));
 sky130_fd_sc_hd__nand2_2 _33389_ (.A(_05168_),
    .B(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__nand2_2 _33390_ (.A(_01040_),
    .B(_03345_),
    .Y(_05171_));
 sky130_fd_sc_hd__xnor2_2 _33391_ (.A(_05170_),
    .B(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__nor2_2 _33392_ (.A(_16257_),
    .B(_18443_),
    .Y(_05173_));
 sky130_fd_sc_hd__and2_2 _33393_ (.A(_04842_),
    .B(_05173_),
    .X(_05175_));
 sky130_fd_sc_hd__a2bb2o_2 _33394_ (.A1_N(_16258_),
    .A2_N(_18200_),
    .B1(_18463_),
    .B2(_16934_),
    .X(_05176_));
 sky130_fd_sc_hd__and2b_2 _33395_ (.A_N(_05175_),
    .B(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__nor2_2 _33396_ (.A(_16619_),
    .B(_04501_),
    .Y(_05178_));
 sky130_fd_sc_hd__xnor2_2 _33397_ (.A(_05177_),
    .B(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__a22o_2 _33398_ (.A1(_04500_),
    .A2(_04842_),
    .B1(_04843_),
    .B2(_04844_),
    .X(_05180_));
 sky130_fd_sc_hd__or2b_2 _33399_ (.A(_05179_),
    .B_N(_05180_),
    .X(_05181_));
 sky130_fd_sc_hd__or2b_2 _33400_ (.A(_05180_),
    .B_N(_05179_),
    .X(_05182_));
 sky130_fd_sc_hd__nand2_2 _33401_ (.A(_05181_),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__xor2_2 _33402_ (.A(_05172_),
    .B(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__a21bo_2 _33403_ (.A1(_04860_),
    .A2(_04863_),
    .B1_N(_04859_),
    .X(_05186_));
 sky130_fd_sc_hd__or4_2 _33404_ (.A(_15173_),
    .B(_15154_),
    .C(_00271_),
    .D(_00666_),
    .X(_05187_));
 sky130_fd_sc_hd__a22o_2 _33405_ (.A1(_15586_),
    .A2(_01647_),
    .B1(_00268_),
    .B2(_01033_),
    .X(_05188_));
 sky130_fd_sc_hd__nand2_2 _33406_ (.A(_05187_),
    .B(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__nor2_2 _33407_ (.A(_03388_),
    .B(_01066_),
    .Y(_05190_));
 sky130_fd_sc_hd__xor2_2 _33408_ (.A(_05189_),
    .B(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__a2bb2o_2 _33409_ (.A1_N(_04879_),
    .A2_N(_04880_),
    .B1(_04881_),
    .B2(_04882_),
    .X(_05192_));
 sky130_fd_sc_hd__and2b_2 _33410_ (.A_N(_05191_),
    .B(_05192_),
    .X(_05193_));
 sky130_fd_sc_hd__and2b_2 _33411_ (.A_N(_05192_),
    .B(_05191_),
    .X(_05194_));
 sky130_fd_sc_hd__nor2_2 _33412_ (.A(_05193_),
    .B(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__xnor2_2 _33413_ (.A(_05186_),
    .B(_05195_),
    .Y(_05197_));
 sky130_fd_sc_hd__and2b_2 _33414_ (.A_N(_04865_),
    .B(_04857_),
    .X(_05198_));
 sky130_fd_sc_hd__a21oi_2 _33415_ (.A1(_04858_),
    .A2(_04864_),
    .B1(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__nor2_2 _33416_ (.A(_05197_),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__and2_2 _33417_ (.A(_05197_),
    .B(_05199_),
    .X(_05201_));
 sky130_fd_sc_hd__nor2_2 _33418_ (.A(_05200_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__xor2_2 _33419_ (.A(_05184_),
    .B(_05202_),
    .X(_05203_));
 sky130_fd_sc_hd__xnor2_2 _33420_ (.A(_05167_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__o21ai_2 _33421_ (.A1(_04868_),
    .A2(_04871_),
    .B1(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__or3_2 _33422_ (.A(_04868_),
    .B(_04871_),
    .C(_05204_),
    .X(_05206_));
 sky130_fd_sc_hd__and2_2 _33423_ (.A(_05205_),
    .B(_05206_),
    .X(_05208_));
 sky130_fd_sc_hd__nand2_2 _33424_ (.A(_14632_),
    .B(_03064_),
    .Y(_05209_));
 sky130_fd_sc_hd__a2bb2o_2 _33425_ (.A1_N(_00589_),
    .A2_N(_04181_),
    .B1(_04005_),
    .B2(_02626_),
    .X(_05210_));
 sky130_fd_sc_hd__nand2_2 _33426_ (.A(_05209_),
    .B(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__nand2_2 _33427_ (.A(_14344_),
    .B(_03064_),
    .Y(_05212_));
 sky130_fd_sc_hd__o211ai_2 _33428_ (.A1(_04899_),
    .A2(_04903_),
    .B1(_05211_),
    .C1(_05212_),
    .Y(_05213_));
 sky130_fd_sc_hd__or2_2 _33429_ (.A(_05212_),
    .B(_05211_),
    .X(_05214_));
 sky130_fd_sc_hd__o31a_2 _33430_ (.A1(_04899_),
    .A2(_04903_),
    .A3(_05211_),
    .B1(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__and4_2 _33431_ (.A(_04904_),
    .B(_04906_),
    .C(_05213_),
    .D(_05215_),
    .X(_05216_));
 sky130_fd_sc_hd__a22o_2 _33432_ (.A1(_04904_),
    .A2(_04906_),
    .B1(_05213_),
    .B2(_05215_),
    .X(_05217_));
 sky130_fd_sc_hd__or2b_2 _33433_ (.A(_05216_),
    .B_N(_05217_),
    .X(_05219_));
 sky130_fd_sc_hd__or2b_2 _33434_ (.A(_04890_),
    .B_N(_04888_),
    .X(_05220_));
 sky130_fd_sc_hd__o21ai_2 _33435_ (.A1(_04883_),
    .A2(_04891_),
    .B1(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__or3_2 _33436_ (.A(_01605_),
    .B(_02647_),
    .C(_04880_),
    .X(_05222_));
 sky130_fd_sc_hd__nor2_2 _33437_ (.A(_02608_),
    .B(_02647_),
    .Y(_05223_));
 sky130_fd_sc_hd__a21o_2 _33438_ (.A1(_14593_),
    .A2(_03438_),
    .B1(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__nand2_2 _33439_ (.A(_05222_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__or3_2 _33440_ (.A(_01028_),
    .B(_01070_),
    .C(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__buf_1 _33441_ (.A(_01070_),
    .X(_05227_));
 sky130_fd_sc_hd__o21ai_2 _33442_ (.A1(_01028_),
    .A2(_05227_),
    .B1(_05225_),
    .Y(_05228_));
 sky130_fd_sc_hd__nand2_2 _33443_ (.A(_05226_),
    .B(_05228_),
    .Y(_05230_));
 sky130_fd_sc_hd__buf_1 _33444_ (.A(_02391_),
    .X(_05231_));
 sky130_fd_sc_hd__nor2_2 _33445_ (.A(_02613_),
    .B(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__nor2_2 _33446_ (.A(_18791_),
    .B(_02643_),
    .Y(_05233_));
 sky130_fd_sc_hd__or3_2 _33447_ (.A(_14626_),
    .B(_02397_),
    .C(_02398_),
    .X(_05234_));
 sky130_fd_sc_hd__xnor2_2 _33448_ (.A(_05233_),
    .B(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__xnor2_2 _33449_ (.A(_05232_),
    .B(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__o31a_2 _33450_ (.A1(_02613_),
    .A2(_04187_),
    .A3(_04886_),
    .B1(_04884_),
    .X(_05237_));
 sky130_fd_sc_hd__xnor2_2 _33451_ (.A(_05236_),
    .B(_05237_),
    .Y(_05238_));
 sky130_fd_sc_hd__xnor2_2 _33452_ (.A(_05230_),
    .B(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__xnor2_2 _33453_ (.A(_04555_),
    .B(_05239_),
    .Y(_05241_));
 sky130_fd_sc_hd__xnor2_2 _33454_ (.A(_05221_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__xnor2_2 _33455_ (.A(_05219_),
    .B(_05242_),
    .Y(_05243_));
 sky130_fd_sc_hd__nor2_2 _33456_ (.A(_04897_),
    .B(_04907_),
    .Y(_05244_));
 sky130_fd_sc_hd__a21oi_2 _33457_ (.A1(_04896_),
    .A2(_04908_),
    .B1(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__xnor2_2 _33458_ (.A(_05243_),
    .B(_05245_),
    .Y(_05246_));
 sky130_fd_sc_hd__xor2_2 _33459_ (.A(_05208_),
    .B(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__nor2_2 _33460_ (.A(_04909_),
    .B(_04912_),
    .Y(_05248_));
 sky130_fd_sc_hd__a21o_2 _33461_ (.A1(_04876_),
    .A2(_04913_),
    .B1(_05248_),
    .X(_05249_));
 sky130_fd_sc_hd__xor2_2 _33462_ (.A(_05247_),
    .B(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__xor2_2 _33463_ (.A(_05166_),
    .B(_05250_),
    .X(_05252_));
 sky130_fd_sc_hd__and2b_2 _33464_ (.A_N(_04916_),
    .B(_04914_),
    .X(_05253_));
 sky130_fd_sc_hd__a21oi_2 _33465_ (.A1(_04830_),
    .A2(_04917_),
    .B1(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__xnor2_2 _33466_ (.A(_05252_),
    .B(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__xnor2_2 _33467_ (.A(_05118_),
    .B(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hd__or2b_2 _33468_ (.A(_04918_),
    .B_N(_04920_),
    .X(_05257_));
 sky130_fd_sc_hd__a21boi_2 _33469_ (.A1(_04776_),
    .A2(_04921_),
    .B1_N(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__xor2_2 _33470_ (.A(_05256_),
    .B(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__xnor2_2 _33471_ (.A(_04774_),
    .B(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__xnor2_2 _33472_ (.A(_05112_),
    .B(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__nand3_2 _33473_ (.A(_05109_),
    .B(_05110_),
    .C(_05261_),
    .Y(_05263_));
 sky130_fd_sc_hd__a21o_2 _33474_ (.A1(_05109_),
    .A2(_05110_),
    .B1(_05261_),
    .X(_05264_));
 sky130_fd_sc_hd__or2b_2 _33475_ (.A(_05079_),
    .B_N(_05080_),
    .X(_05265_));
 sky130_fd_sc_hd__and2b_2 _33476_ (.A_N(_05000_),
    .B(_04998_),
    .X(_05266_));
 sky130_fd_sc_hd__a21oi_2 _33477_ (.A1(_04993_),
    .A2(_05001_),
    .B1(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__and4_2 _33478_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[58]),
    .D(iX[59]),
    .X(_05268_));
 sky130_fd_sc_hd__a22oi_2 _33479_ (.A1(iY[45]),
    .A2(iX[58]),
    .B1(iX[59]),
    .B2(iY[44]),
    .Y(_05269_));
 sky130_fd_sc_hd__nor2_2 _33480_ (.A(_05268_),
    .B(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__nand2_2 _33481_ (.A(iY[46]),
    .B(iX[57]),
    .Y(_05271_));
 sky130_fd_sc_hd__xnor2_2 _33482_ (.A(_05270_),
    .B(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__and2_2 _33483_ (.A(iY[42]),
    .B(iX[62]),
    .X(_05274_));
 sky130_fd_sc_hd__nand3_2 _33484_ (.A(iY[41]),
    .B(iX[61]),
    .C(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__a22o_2 _33485_ (.A1(iY[42]),
    .A2(iX[61]),
    .B1(iX[62]),
    .B2(iY[41]),
    .X(_05276_));
 sky130_fd_sc_hd__and2_2 _33486_ (.A(iY[43]),
    .B(iX[60]),
    .X(_05277_));
 sky130_fd_sc_hd__a21oi_2 _33487_ (.A1(_05275_),
    .A2(_05276_),
    .B1(_05277_),
    .Y(_05278_));
 sky130_fd_sc_hd__and3_2 _33488_ (.A(_05275_),
    .B(_05276_),
    .C(_05277_),
    .X(_05279_));
 sky130_fd_sc_hd__nor2_2 _33489_ (.A(_05278_),
    .B(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__o21ba_2 _33490_ (.A1(_04995_),
    .A2(_04997_),
    .B1_N(_04994_),
    .X(_05281_));
 sky130_fd_sc_hd__xnor2_2 _33491_ (.A(_05280_),
    .B(_05281_),
    .Y(_05282_));
 sky130_fd_sc_hd__xnor2_2 _33492_ (.A(_05272_),
    .B(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__or2_2 _33493_ (.A(_04984_),
    .B(_05283_),
    .X(_05285_));
 sky130_fd_sc_hd__nand2_2 _33494_ (.A(_04984_),
    .B(_05283_),
    .Y(_05286_));
 sky130_fd_sc_hd__and2_2 _33495_ (.A(_05285_),
    .B(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__xnor2_2 _33496_ (.A(_05267_),
    .B(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__or3b_2 _33497_ (.A(_04596_),
    .B(_04980_),
    .C_N(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__a31o_2 _33498_ (.A1(iY[40]),
    .A2(iX[63]),
    .A3(_04239_),
    .B1(_05288_),
    .X(_05290_));
 sky130_fd_sc_hd__nand2_2 _33499_ (.A(_05289_),
    .B(_05290_),
    .Y(_05291_));
 sky130_fd_sc_hd__xnor2_2 _33500_ (.A(_05008_),
    .B(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__inv_2 _33501_ (.A(_04970_),
    .Y(_05293_));
 sky130_fd_sc_hd__and4_2 _33502_ (.A(iX[49]),
    .B(iX[50]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_05294_));
 sky130_fd_sc_hd__a22oi_2 _33503_ (.A1(iX[50]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[49]),
    .Y(_05296_));
 sky130_fd_sc_hd__nor2_2 _33504_ (.A(_05294_),
    .B(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__nand2_2 _33505_ (.A(iX[48]),
    .B(iY[55]),
    .Y(_05298_));
 sky130_fd_sc_hd__xnor2_2 _33506_ (.A(_05297_),
    .B(_05298_),
    .Y(_05299_));
 sky130_fd_sc_hd__and4_2 _33507_ (.A(iY[50]),
    .B(iY[51]),
    .C(iX[52]),
    .D(iX[53]),
    .X(_05300_));
 sky130_fd_sc_hd__a22oi_2 _33508_ (.A1(iY[51]),
    .A2(iX[52]),
    .B1(iX[53]),
    .B2(iY[50]),
    .Y(_05301_));
 sky130_fd_sc_hd__nor2_2 _33509_ (.A(_05300_),
    .B(_05301_),
    .Y(_05302_));
 sky130_fd_sc_hd__nand2_2 _33510_ (.A(iX[51]),
    .B(iY[52]),
    .Y(_05303_));
 sky130_fd_sc_hd__xnor2_2 _33511_ (.A(_05302_),
    .B(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__o21ba_2 _33512_ (.A1(_04947_),
    .A2(_04949_),
    .B1_N(_04946_),
    .X(_05305_));
 sky130_fd_sc_hd__xnor2_2 _33513_ (.A(_05304_),
    .B(_05305_),
    .Y(_05307_));
 sky130_fd_sc_hd__and2_2 _33514_ (.A(_05299_),
    .B(_05307_),
    .X(_05308_));
 sky130_fd_sc_hd__nor2_2 _33515_ (.A(_05299_),
    .B(_05307_),
    .Y(_05309_));
 sky130_fd_sc_hd__or2_2 _33516_ (.A(_05308_),
    .B(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__or3_2 _33517_ (.A(_04958_),
    .B(_04962_),
    .C(_04963_),
    .X(_05311_));
 sky130_fd_sc_hd__o21ba_2 _33518_ (.A1(_04990_),
    .A2(_04992_),
    .B1_N(_04989_),
    .X(_05312_));
 sky130_fd_sc_hd__and4_2 _33519_ (.A(iY[47]),
    .B(iY[48]),
    .C(iX[55]),
    .D(iX[56]),
    .X(_05313_));
 sky130_fd_sc_hd__a22oi_2 _33520_ (.A1(iY[48]),
    .A2(iX[55]),
    .B1(iX[56]),
    .B2(iY[47]),
    .Y(_05314_));
 sky130_fd_sc_hd__nand2_2 _33521_ (.A(iY[49]),
    .B(iX[54]),
    .Y(_05315_));
 sky130_fd_sc_hd__o21a_2 _33522_ (.A1(_05313_),
    .A2(_05314_),
    .B1(_05315_),
    .X(_05316_));
 sky130_fd_sc_hd__nor3_2 _33523_ (.A(_05313_),
    .B(_05314_),
    .C(_05315_),
    .Y(_05318_));
 sky130_fd_sc_hd__nor2_2 _33524_ (.A(_05316_),
    .B(_05318_),
    .Y(_05319_));
 sky130_fd_sc_hd__xnor2_2 _33525_ (.A(_05312_),
    .B(_05319_),
    .Y(_05320_));
 sky130_fd_sc_hd__o21ai_2 _33526_ (.A1(_04959_),
    .A2(_04963_),
    .B1(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__or3_2 _33527_ (.A(_04959_),
    .B(_04963_),
    .C(_05320_),
    .X(_05322_));
 sky130_fd_sc_hd__nand2_2 _33528_ (.A(_05321_),
    .B(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__a21oi_2 _33529_ (.A1(_05311_),
    .A2(_04967_),
    .B1(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__and3_2 _33530_ (.A(_05311_),
    .B(_04967_),
    .C(_05323_),
    .X(_05325_));
 sky130_fd_sc_hd__or3_2 _33531_ (.A(_05310_),
    .B(_05324_),
    .C(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__o21ai_2 _33532_ (.A1(_05324_),
    .A2(_05325_),
    .B1(_05310_),
    .Y(_05327_));
 sky130_fd_sc_hd__nand2_2 _33533_ (.A(_05326_),
    .B(_05327_),
    .Y(_05329_));
 sky130_fd_sc_hd__a21oi_2 _33534_ (.A1(_05003_),
    .A2(_05006_),
    .B1(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__and3_2 _33535_ (.A(_05003_),
    .B(_05006_),
    .C(_05329_),
    .X(_05331_));
 sky130_fd_sc_hd__a211o_2 _33536_ (.A1(_05293_),
    .A2(_04972_),
    .B1(_05330_),
    .C1(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__o211ai_2 _33537_ (.A1(_05330_),
    .A2(_05331_),
    .B1(_05293_),
    .C1(_04972_),
    .Y(_05333_));
 sky130_fd_sc_hd__nand3_2 _33538_ (.A(_05292_),
    .B(_05332_),
    .C(_05333_),
    .Y(_05334_));
 sky130_fd_sc_hd__a21o_2 _33539_ (.A1(_05332_),
    .A2(_05333_),
    .B1(_05292_),
    .X(_05335_));
 sky130_fd_sc_hd__nand2_2 _33540_ (.A(_05334_),
    .B(_05335_),
    .Y(_05336_));
 sky130_fd_sc_hd__a21oi_2 _33541_ (.A1(_05011_),
    .A2(_05015_),
    .B1(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__and3_2 _33542_ (.A(_05011_),
    .B(_05015_),
    .C(_05336_),
    .X(_05338_));
 sky130_fd_sc_hd__inv_2 _33543_ (.A(_05058_),
    .Y(_05340_));
 sky130_fd_sc_hd__or2b_2 _33544_ (.A(_05027_),
    .B_N(_05026_),
    .X(_05341_));
 sky130_fd_sc_hd__and4_2 _33545_ (.A(iX[43]),
    .B(iX[44]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_05342_));
 sky130_fd_sc_hd__a22oi_2 _33546_ (.A1(iX[44]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[43]),
    .Y(_05343_));
 sky130_fd_sc_hd__nor2_2 _33547_ (.A(_05342_),
    .B(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__nand2_2 _33548_ (.A(iX[42]),
    .B(iY[61]),
    .Y(_05345_));
 sky130_fd_sc_hd__xnor2_2 _33549_ (.A(_05344_),
    .B(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__o21ba_2 _33550_ (.A1(_05023_),
    .A2(_05025_),
    .B1_N(_05022_),
    .X(_05347_));
 sky130_fd_sc_hd__xnor2_2 _33551_ (.A(_05346_),
    .B(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__nand2_2 _33552_ (.A(iX[41]),
    .B(iY[62]),
    .Y(_05349_));
 sky130_fd_sc_hd__xor2_2 _33553_ (.A(_05348_),
    .B(_05349_),
    .X(_05351_));
 sky130_fd_sc_hd__a21oi_2 _33554_ (.A1(_05341_),
    .A2(_05031_),
    .B1(_05351_),
    .Y(_05352_));
 sky130_fd_sc_hd__and3_2 _33555_ (.A(_05341_),
    .B(_05031_),
    .C(_05351_),
    .X(_05353_));
 sky130_fd_sc_hd__nor2_2 _33556_ (.A(_05352_),
    .B(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__nand2_2 _33557_ (.A(iX[40]),
    .B(iY[63]),
    .Y(_05355_));
 sky130_fd_sc_hd__xnor2_2 _33558_ (.A(_05354_),
    .B(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__or2b_2 _33559_ (.A(_05044_),
    .B_N(_05049_),
    .X(_05357_));
 sky130_fd_sc_hd__or2b_2 _33560_ (.A(_05042_),
    .B_N(_05050_),
    .X(_05358_));
 sky130_fd_sc_hd__and2b_2 _33561_ (.A_N(_04951_),
    .B(_04950_),
    .X(_05359_));
 sky130_fd_sc_hd__o21ba_2 _33562_ (.A1(_05046_),
    .A2(_05048_),
    .B1_N(_05045_),
    .X(_05360_));
 sky130_fd_sc_hd__o21ba_2 _33563_ (.A1(_04941_),
    .A2(_04943_),
    .B1_N(_04940_),
    .X(_05362_));
 sky130_fd_sc_hd__and4_2 _33564_ (.A(iX[46]),
    .B(iX[47]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_05363_));
 sky130_fd_sc_hd__a22oi_2 _33565_ (.A1(iX[47]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[46]),
    .Y(_05364_));
 sky130_fd_sc_hd__nor2_2 _33566_ (.A(_05363_),
    .B(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__nand2_2 _33567_ (.A(iX[45]),
    .B(iY[58]),
    .Y(_05366_));
 sky130_fd_sc_hd__xnor2_2 _33568_ (.A(_05365_),
    .B(_05366_),
    .Y(_05367_));
 sky130_fd_sc_hd__xnor2_2 _33569_ (.A(_05362_),
    .B(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__xnor2_2 _33570_ (.A(_05360_),
    .B(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__o21a_2 _33571_ (.A1(_05359_),
    .A2(_04953_),
    .B1(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__nor3_2 _33572_ (.A(_05359_),
    .B(_04953_),
    .C(_05369_),
    .Y(_05371_));
 sky130_fd_sc_hd__a211oi_2 _33573_ (.A1(_05357_),
    .A2(_05358_),
    .B1(_05370_),
    .C1(_05371_),
    .Y(_05373_));
 sky130_fd_sc_hd__o211a_2 _33574_ (.A1(_05370_),
    .A2(_05371_),
    .B1(_05357_),
    .C1(_05358_),
    .X(_05374_));
 sky130_fd_sc_hd__nor2_2 _33575_ (.A(_05052_),
    .B(_05055_),
    .Y(_05375_));
 sky130_fd_sc_hd__or3_2 _33576_ (.A(_05373_),
    .B(_05374_),
    .C(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__o21ai_2 _33577_ (.A1(_05373_),
    .A2(_05374_),
    .B1(_05375_),
    .Y(_05377_));
 sky130_fd_sc_hd__and3_2 _33578_ (.A(_05356_),
    .B(_05376_),
    .C(_05377_),
    .X(_05378_));
 sky130_fd_sc_hd__a21oi_2 _33579_ (.A1(_05376_),
    .A2(_05377_),
    .B1(_05356_),
    .Y(_05379_));
 sky130_fd_sc_hd__nor2_2 _33580_ (.A(_05378_),
    .B(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__o21ai_2 _33581_ (.A1(_04975_),
    .A2(_04978_),
    .B1(_05380_),
    .Y(_05381_));
 sky130_fd_sc_hd__or3_2 _33582_ (.A(_04975_),
    .B(_04978_),
    .C(_05380_),
    .X(_05382_));
 sky130_fd_sc_hd__o211ai_2 _33583_ (.A1(_05340_),
    .A2(_05060_),
    .B1(_05381_),
    .C1(_05382_),
    .Y(_05384_));
 sky130_fd_sc_hd__a211o_2 _33584_ (.A1(_05381_),
    .A2(_05382_),
    .B1(_05340_),
    .C1(_05060_),
    .X(_05385_));
 sky130_fd_sc_hd__or4bb_2 _33585_ (.A(_05337_),
    .B(_05338_),
    .C_N(_05384_),
    .D_N(_05385_),
    .X(_05386_));
 sky130_fd_sc_hd__a2bb2o_2 _33586_ (.A1_N(_05337_),
    .A2_N(_05338_),
    .B1(_05384_),
    .B2(_05385_),
    .X(_05387_));
 sky130_fd_sc_hd__a21bo_2 _33587_ (.A1(_05016_),
    .A2(_05017_),
    .B1_N(_05068_),
    .X(_05388_));
 sky130_fd_sc_hd__and3_2 _33588_ (.A(_05386_),
    .B(_05387_),
    .C(_05388_),
    .X(_05389_));
 sky130_fd_sc_hd__a21oi_2 _33589_ (.A1(_05386_),
    .A2(_05387_),
    .B1(_05388_),
    .Y(_05390_));
 sky130_fd_sc_hd__or2_2 _33590_ (.A(_05389_),
    .B(_05390_),
    .X(_05391_));
 sky130_fd_sc_hd__o21ai_2 _33591_ (.A1(_05019_),
    .A2(_05066_),
    .B1(_05063_),
    .Y(_05392_));
 sky130_fd_sc_hd__xnor2_2 _33592_ (.A(_05391_),
    .B(_05392_),
    .Y(_05393_));
 sky130_fd_sc_hd__and2b_2 _33593_ (.A_N(_05073_),
    .B(_05074_),
    .X(_05395_));
 sky130_fd_sc_hd__o21ba_2 _33594_ (.A1(_05070_),
    .A2(_05072_),
    .B1_N(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__xor2_2 _33595_ (.A(_05393_),
    .B(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__a31o_2 _33596_ (.A1(iX[39]),
    .A2(iY[63]),
    .A3(_05036_),
    .B1(_05034_),
    .X(_05398_));
 sky130_fd_sc_hd__xor2_2 _33597_ (.A(_05397_),
    .B(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__nand3_2 _33598_ (.A(_05077_),
    .B(_05265_),
    .C(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__a21oi_2 _33599_ (.A1(_05077_),
    .A2(_05265_),
    .B1(_05399_),
    .Y(_05401_));
 sky130_fd_sc_hd__inv_2 _33600_ (.A(_05401_),
    .Y(_05402_));
 sky130_fd_sc_hd__nand2_2 _33601_ (.A(_05400_),
    .B(_05402_),
    .Y(_05403_));
 sky130_fd_sc_hd__a21oi_2 _33602_ (.A1(_05082_),
    .A2(_05083_),
    .B1(_05081_),
    .Y(_05404_));
 sky130_fd_sc_hd__o21ba_2 _33603_ (.A1(_05085_),
    .A2(_05089_),
    .B1_N(_05404_),
    .X(_05406_));
 sky130_fd_sc_hd__xnor2_2 _33604_ (.A(_05403_),
    .B(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__a21o_2 _33605_ (.A1(_05263_),
    .A2(_05264_),
    .B1(_05407_),
    .X(_05408_));
 sky130_fd_sc_hd__nand3_2 _33606_ (.A(_05263_),
    .B(_05264_),
    .C(_05407_),
    .Y(_05409_));
 sky130_fd_sc_hd__nand3_2 _33607_ (.A(_13064_),
    .B(_05408_),
    .C(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__a21o_2 _33608_ (.A1(_05408_),
    .A2(_05409_),
    .B1(_13064_),
    .X(_05411_));
 sky130_fd_sc_hd__nor2_2 _33609_ (.A(_04937_),
    .B(_05090_),
    .Y(_05412_));
 sky130_fd_sc_hd__a21o_2 _33610_ (.A1(_04769_),
    .A2(_05092_),
    .B1(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__a21o_2 _33611_ (.A1(_05410_),
    .A2(_05411_),
    .B1(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__nand3_2 _33612_ (.A(_05413_),
    .B(_05410_),
    .C(_05411_),
    .Y(_05415_));
 sky130_fd_sc_hd__nand2_2 _33613_ (.A(_05414_),
    .B(_05415_),
    .Y(_05417_));
 sky130_fd_sc_hd__xnor2_2 _33614_ (.A(_05107_),
    .B(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__xor2_2 _33615_ (.A(_12911_),
    .B(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__o21ai_2 _33616_ (.A1(_05102_),
    .A2(_05105_),
    .B1(_05100_),
    .Y(_05420_));
 sky130_fd_sc_hd__xnor2_2 _33617_ (.A(_05419_),
    .B(_05420_),
    .Y(oO[71]));
 sky130_fd_sc_hd__a2111o_2 _33618_ (.A1(_04055_),
    .A2(_04059_),
    .B1(_04930_),
    .C1(_04931_),
    .D1(_05261_),
    .X(_05421_));
 sky130_fd_sc_hd__nor2_2 _33619_ (.A(_05112_),
    .B(_05260_),
    .Y(_05422_));
 sky130_fd_sc_hd__or3_2 _33620_ (.A(_04930_),
    .B(_04935_),
    .C(_05261_),
    .X(_05423_));
 sky130_fd_sc_hd__a21o_2 _33621_ (.A1(_05112_),
    .A2(_05260_),
    .B1(_05109_),
    .X(_05424_));
 sky130_fd_sc_hd__and3b_2 _33622_ (.A_N(_05422_),
    .B(_05423_),
    .C(_05424_),
    .X(_05425_));
 sky130_fd_sc_hd__and2b_2 _33623_ (.A_N(_05122_),
    .B(_05164_),
    .X(_05427_));
 sky130_fd_sc_hd__and2b_2 _33624_ (.A_N(_05121_),
    .B(_05165_),
    .X(_05428_));
 sky130_fd_sc_hd__or2_2 _33625_ (.A(_05427_),
    .B(_05428_),
    .X(_05429_));
 sky130_fd_sc_hd__and3_2 _33626_ (.A(_05136_),
    .B(_05137_),
    .C(_05139_),
    .X(_05430_));
 sky130_fd_sc_hd__and2_2 _33627_ (.A(_05123_),
    .B(_05140_),
    .X(_05431_));
 sky130_fd_sc_hd__nor2_2 _33628_ (.A(_05430_),
    .B(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__xnor2_2 _33629_ (.A(_05429_),
    .B(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__and2b_2 _33630_ (.A_N(_05159_),
    .B(_05161_),
    .X(_05434_));
 sky130_fd_sc_hd__or3_2 _33631_ (.A(_05157_),
    .B(_05158_),
    .C(_05161_),
    .X(_05435_));
 sky130_fd_sc_hd__o21ai_2 _33632_ (.A1(_05142_),
    .A2(_05434_),
    .B1(_05435_),
    .Y(_05436_));
 sky130_fd_sc_hd__or2b_2 _33633_ (.A(_05167_),
    .B_N(_05203_),
    .X(_05438_));
 sky130_fd_sc_hd__nand2_2 _33634_ (.A(_05438_),
    .B(_05205_),
    .Y(_05439_));
 sky130_fd_sc_hd__buf_1 _33635_ (.A(_03318_),
    .X(_05440_));
 sky130_fd_sc_hd__buf_1 _33636_ (.A(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__or2_2 _33637_ (.A(_04785_),
    .B(_05124_),
    .X(_05442_));
 sky130_fd_sc_hd__o31a_2 _33638_ (.A1(_00990_),
    .A2(_05441_),
    .A3(_05125_),
    .B1(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__or3_2 _33639_ (.A(_01576_),
    .B(_02317_),
    .C(_05124_),
    .X(_05444_));
 sky130_fd_sc_hd__a2bb2o_2 _33640_ (.A1_N(_01797_),
    .A2_N(_02317_),
    .B1(_02928_),
    .B2(_18157_),
    .X(_05445_));
 sky130_fd_sc_hd__nand2_2 _33641_ (.A(_05444_),
    .B(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__nor2_2 _33642_ (.A(_16288_),
    .B(_03318_),
    .Y(_05447_));
 sky130_fd_sc_hd__xnor2_2 _33643_ (.A(_05446_),
    .B(_05447_),
    .Y(_05449_));
 sky130_fd_sc_hd__buf_1 _33644_ (.A(_01757_),
    .X(_05450_));
 sky130_fd_sc_hd__nand2_2 _33645_ (.A(_02983_),
    .B(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__nand2_2 _33646_ (.A(_02994_),
    .B(_00566_),
    .Y(_05452_));
 sky130_fd_sc_hd__a22o_2 _33647_ (.A1(_02994_),
    .A2(_05450_),
    .B1(_00566_),
    .B2(_02983_),
    .X(_05453_));
 sky130_fd_sc_hd__o21ai_2 _33648_ (.A1(_05451_),
    .A2(_05452_),
    .B1(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__nand2_2 _33649_ (.A(_15888_),
    .B(_03327_),
    .Y(_05455_));
 sky130_fd_sc_hd__xnor2_2 _33650_ (.A(_05454_),
    .B(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__o21a_2 _33651_ (.A1(_05131_),
    .A2(_05132_),
    .B1(_05128_),
    .X(_05457_));
 sky130_fd_sc_hd__nor2_2 _33652_ (.A(_05456_),
    .B(_05457_),
    .Y(_05458_));
 sky130_fd_sc_hd__nand2_2 _33653_ (.A(_05456_),
    .B(_05457_),
    .Y(_05460_));
 sky130_fd_sc_hd__and2b_2 _33654_ (.A_N(_05458_),
    .B(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__xnor2_2 _33655_ (.A(_05449_),
    .B(_05461_),
    .Y(_05462_));
 sky130_fd_sc_hd__o21ai_2 _33656_ (.A1(_05133_),
    .A2(_05134_),
    .B1(_05136_),
    .Y(_05463_));
 sky130_fd_sc_hd__xnor2_2 _33657_ (.A(_05462_),
    .B(_05463_),
    .Y(_05464_));
 sky130_fd_sc_hd__xnor2_2 _33658_ (.A(_05443_),
    .B(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__and2_2 _33659_ (.A(_05146_),
    .B(_05155_),
    .X(_05466_));
 sky130_fd_sc_hd__or2b_2 _33660_ (.A(_05153_),
    .B_N(_05148_),
    .X(_05467_));
 sky130_fd_sc_hd__or2b_2 _33661_ (.A(_05154_),
    .B_N(_05147_),
    .X(_05468_));
 sky130_fd_sc_hd__nand2_2 _33662_ (.A(_05467_),
    .B(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__o21ai_2 _33663_ (.A1(_05172_),
    .A2(_05183_),
    .B1(_05181_),
    .Y(_05471_));
 sky130_fd_sc_hd__or3b_2 _33664_ (.A(_02471_),
    .B(_03341_),
    .C_N(_05150_),
    .X(_05472_));
 sky130_fd_sc_hd__o21ai_2 _33665_ (.A1(_04813_),
    .A2(_05149_),
    .B1(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__o21ai_2 _33666_ (.A1(_05170_),
    .A2(_05171_),
    .B1(_05168_),
    .Y(_05474_));
 sky130_fd_sc_hd__nand2_2 _33667_ (.A(_00633_),
    .B(_18734_),
    .Y(_05475_));
 sky130_fd_sc_hd__or3_2 _33668_ (.A(_01828_),
    .B(_18111_),
    .C(_18113_),
    .X(_05476_));
 sky130_fd_sc_hd__xor2_2 _33669_ (.A(_05475_),
    .B(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__nor2_2 _33670_ (.A(_03378_),
    .B(_03341_),
    .Y(_05478_));
 sky130_fd_sc_hd__xnor2_2 _33671_ (.A(_05477_),
    .B(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__xnor2_2 _33672_ (.A(_05474_),
    .B(_05479_),
    .Y(_05480_));
 sky130_fd_sc_hd__xnor2_2 _33673_ (.A(_05473_),
    .B(_05480_),
    .Y(_05482_));
 sky130_fd_sc_hd__xor2_2 _33674_ (.A(_05471_),
    .B(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__xnor2_2 _33675_ (.A(_05469_),
    .B(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__o21a_2 _33676_ (.A1(_05466_),
    .A2(_05157_),
    .B1(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__nor3_2 _33677_ (.A(_05466_),
    .B(_05157_),
    .C(_05484_),
    .Y(_05486_));
 sky130_fd_sc_hd__nor2_2 _33678_ (.A(_05485_),
    .B(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__xnor2_2 _33679_ (.A(_05465_),
    .B(_05487_),
    .Y(_05488_));
 sky130_fd_sc_hd__xor2_2 _33680_ (.A(_05439_),
    .B(_05488_),
    .X(_05489_));
 sky130_fd_sc_hd__xor2_2 _33681_ (.A(_05436_),
    .B(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__a21oi_2 _33682_ (.A1(_05184_),
    .A2(_05202_),
    .B1(_05200_),
    .Y(_05491_));
 sky130_fd_sc_hd__or2b_2 _33683_ (.A(_05241_),
    .B_N(_05221_),
    .X(_05493_));
 sky130_fd_sc_hd__o21ai_2 _33684_ (.A1(_04555_),
    .A2(_05239_),
    .B1(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__or2_2 _33685_ (.A(_18363_),
    .B(_01058_),
    .X(_05495_));
 sky130_fd_sc_hd__or3_2 _33686_ (.A(_00649_),
    .B(_17409_),
    .C(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__o21ai_2 _33687_ (.A1(_00649_),
    .A2(_17409_),
    .B1(_05495_),
    .Y(_05497_));
 sky130_fd_sc_hd__and2_2 _33688_ (.A(_05496_),
    .B(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__a21o_2 _33689_ (.A1(_04837_),
    .A2(_03345_),
    .B1(_05498_),
    .X(_05499_));
 sky130_fd_sc_hd__buf_1 _33690_ (.A(_17628_),
    .X(_05500_));
 sky130_fd_sc_hd__or3b_2 _33691_ (.A(_04504_),
    .B(_05500_),
    .C_N(_05498_),
    .X(_05501_));
 sky130_fd_sc_hd__nand2_2 _33692_ (.A(_05499_),
    .B(_05501_),
    .Y(_05502_));
 sky130_fd_sc_hd__buf_1 _33693_ (.A(_01066_),
    .X(_05504_));
 sky130_fd_sc_hd__nor2_2 _33694_ (.A(_01804_),
    .B(_05504_),
    .Y(_05505_));
 sky130_fd_sc_hd__xnor2_2 _33695_ (.A(_05173_),
    .B(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__buf_1 _33696_ (.A(_18209_),
    .X(_05507_));
 sky130_fd_sc_hd__nand2_2 _33697_ (.A(_16614_),
    .B(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__xnor2_2 _33698_ (.A(_05506_),
    .B(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__a21o_2 _33699_ (.A1(_05176_),
    .A2(_05178_),
    .B1(_05175_),
    .X(_05510_));
 sky130_fd_sc_hd__or2b_2 _33700_ (.A(_05509_),
    .B_N(_05510_),
    .X(_05511_));
 sky130_fd_sc_hd__or2b_2 _33701_ (.A(_05510_),
    .B_N(_05509_),
    .X(_05512_));
 sky130_fd_sc_hd__nand2_2 _33702_ (.A(_05511_),
    .B(_05512_),
    .Y(_05513_));
 sky130_fd_sc_hd__xor2_2 _33703_ (.A(_05502_),
    .B(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__a21bo_2 _33704_ (.A1(_05188_),
    .A2(_05190_),
    .B1_N(_05187_),
    .X(_05515_));
 sky130_fd_sc_hd__nand2_2 _33705_ (.A(_05222_),
    .B(_05226_),
    .Y(_05516_));
 sky130_fd_sc_hd__nand2_2 _33706_ (.A(_15586_),
    .B(_02629_),
    .Y(_05517_));
 sky130_fd_sc_hd__or3_2 _33707_ (.A(_14949_),
    .B(_04162_),
    .C(_05517_),
    .X(_05518_));
 sky130_fd_sc_hd__a22o_2 _33708_ (.A1(_15586_),
    .A2(_01862_),
    .B1(_02629_),
    .B2(_01033_),
    .X(_05519_));
 sky130_fd_sc_hd__nand2_2 _33709_ (.A(_05518_),
    .B(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__buf_1 _33710_ (.A(_03388_),
    .X(_05521_));
 sky130_fd_sc_hd__buf_1 _33711_ (.A(_00271_),
    .X(_05522_));
 sky130_fd_sc_hd__nor2_2 _33712_ (.A(_05521_),
    .B(_05522_),
    .Y(_05523_));
 sky130_fd_sc_hd__xor2_2 _33713_ (.A(_05520_),
    .B(_05523_),
    .X(_05525_));
 sky130_fd_sc_hd__xnor2_2 _33714_ (.A(_05516_),
    .B(_05525_),
    .Y(_05526_));
 sky130_fd_sc_hd__xnor2_2 _33715_ (.A(_05515_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__a21oi_2 _33716_ (.A1(_05186_),
    .A2(_05195_),
    .B1(_05193_),
    .Y(_05528_));
 sky130_fd_sc_hd__xor2_2 _33717_ (.A(_05527_),
    .B(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__xnor2_2 _33718_ (.A(_05514_),
    .B(_05529_),
    .Y(_05530_));
 sky130_fd_sc_hd__xnor2_2 _33719_ (.A(_05494_),
    .B(_05530_),
    .Y(_05531_));
 sky130_fd_sc_hd__xnor2_2 _33720_ (.A(_05491_),
    .B(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__buf_1 _33721_ (.A(_03064_),
    .X(_05533_));
 sky130_fd_sc_hd__o22a_2 _33722_ (.A1(_00990_),
    .A2(_04181_),
    .B1(_04901_),
    .B2(_14626_),
    .X(_05534_));
 sky130_fd_sc_hd__a21o_2 _33723_ (.A1(_15641_),
    .A2(_05533_),
    .B1(_05534_),
    .X(_05536_));
 sky130_fd_sc_hd__a21o_2 _33724_ (.A1(_05209_),
    .A2(_05215_),
    .B1(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__nand3_2 _33725_ (.A(_05209_),
    .B(_05215_),
    .C(_05536_),
    .Y(_05538_));
 sky130_fd_sc_hd__and3_2 _33726_ (.A(_14593_),
    .B(_03994_),
    .C(_05223_),
    .X(_05539_));
 sky130_fd_sc_hd__o22a_2 _33727_ (.A1(_01605_),
    .A2(_02647_),
    .B1(_02391_),
    .B2(_02608_),
    .X(_05540_));
 sky130_fd_sc_hd__or2_2 _33728_ (.A(_05539_),
    .B(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__and3b_2 _33729_ (.A_N(_05541_),
    .B(_03438_),
    .C(_03023_),
    .X(_05542_));
 sky130_fd_sc_hd__buf_1 _33730_ (.A(_01866_),
    .X(_05543_));
 sky130_fd_sc_hd__o21a_2 _33731_ (.A1(_01028_),
    .A2(_05543_),
    .B1(_05541_),
    .X(_05544_));
 sky130_fd_sc_hd__nor2_2 _33732_ (.A(_05542_),
    .B(_05544_),
    .Y(_05545_));
 sky130_fd_sc_hd__inv_2 _33733_ (.A(_05233_),
    .Y(_05547_));
 sky130_fd_sc_hd__or2_2 _33734_ (.A(_05547_),
    .B(_05234_),
    .X(_05548_));
 sky130_fd_sc_hd__a21boi_2 _33735_ (.A1(_05232_),
    .A2(_05235_),
    .B1_N(_05548_),
    .Y(_05549_));
 sky130_fd_sc_hd__buf_1 _33736_ (.A(_02652_),
    .X(_05550_));
 sky130_fd_sc_hd__a22o_2 _33737_ (.A1(_13889_),
    .A2(_03458_),
    .B1(_03454_),
    .B2(_13544_),
    .X(_05551_));
 sky130_fd_sc_hd__o31a_2 _33738_ (.A1(_02613_),
    .A2(_05550_),
    .A3(_05547_),
    .B1(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__and2b_2 _33739_ (.A_N(_05549_),
    .B(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__and2b_2 _33740_ (.A_N(_05552_),
    .B(_05549_),
    .X(_05554_));
 sky130_fd_sc_hd__nor2_2 _33741_ (.A(_05553_),
    .B(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__xnor2_2 _33742_ (.A(_05545_),
    .B(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hd__or2_2 _33743_ (.A(_05236_),
    .B(_05237_),
    .X(_05558_));
 sky130_fd_sc_hd__o21ai_2 _33744_ (.A1(_05230_),
    .A2(_05238_),
    .B1(_05558_),
    .Y(_05559_));
 sky130_fd_sc_hd__xnor2_2 _33745_ (.A(_05556_),
    .B(_05559_),
    .Y(_05560_));
 sky130_fd_sc_hd__nand3_2 _33746_ (.A(_05537_),
    .B(_05538_),
    .C(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__a21o_2 _33747_ (.A1(_05537_),
    .A2(_05538_),
    .B1(_05560_),
    .X(_05562_));
 sky130_fd_sc_hd__a21o_2 _33748_ (.A1(_05217_),
    .A2(_05242_),
    .B1(_05216_),
    .X(_05563_));
 sky130_fd_sc_hd__and3_2 _33749_ (.A(_05561_),
    .B(_05562_),
    .C(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__a21oi_2 _33750_ (.A1(_05561_),
    .A2(_05562_),
    .B1(_05563_),
    .Y(_05565_));
 sky130_fd_sc_hd__nor2_2 _33751_ (.A(_05564_),
    .B(_05565_),
    .Y(_05566_));
 sky130_fd_sc_hd__xnor2_2 _33752_ (.A(_05532_),
    .B(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__and2b_2 _33753_ (.A_N(_05245_),
    .B(_05243_),
    .X(_05569_));
 sky130_fd_sc_hd__a21oi_2 _33754_ (.A1(_05208_),
    .A2(_05246_),
    .B1(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__xnor2_2 _33755_ (.A(_05567_),
    .B(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__xor2_2 _33756_ (.A(_05490_),
    .B(_05571_),
    .X(_05572_));
 sky130_fd_sc_hd__nand2_2 _33757_ (.A(_05247_),
    .B(_05249_),
    .Y(_05573_));
 sky130_fd_sc_hd__a21boi_2 _33758_ (.A1(_05166_),
    .A2(_05250_),
    .B1_N(_05573_),
    .Y(_05574_));
 sky130_fd_sc_hd__xnor2_2 _33759_ (.A(_05572_),
    .B(_05574_),
    .Y(_05575_));
 sky130_fd_sc_hd__xnor2_2 _33760_ (.A(_05433_),
    .B(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hd__or2b_2 _33761_ (.A(_05254_),
    .B_N(_05252_),
    .X(_05577_));
 sky130_fd_sc_hd__a21boi_2 _33762_ (.A1(_05118_),
    .A2(_05255_),
    .B1_N(_05577_),
    .Y(_05578_));
 sky130_fd_sc_hd__nor2_2 _33763_ (.A(_05576_),
    .B(_05578_),
    .Y(_05580_));
 sky130_fd_sc_hd__and2_2 _33764_ (.A(_05576_),
    .B(_05578_),
    .X(_05581_));
 sky130_fd_sc_hd__nor2_2 _33765_ (.A(_05580_),
    .B(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__xnor2_2 _33766_ (.A(_05116_),
    .B(_05582_),
    .Y(_05583_));
 sky130_fd_sc_hd__nor2_2 _33767_ (.A(_05256_),
    .B(_05258_),
    .Y(_05584_));
 sky130_fd_sc_hd__a21oi_2 _33768_ (.A1(_04774_),
    .A2(_05259_),
    .B1(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__nor2_2 _33769_ (.A(_05583_),
    .B(_05585_),
    .Y(_05586_));
 sky130_fd_sc_hd__and2_2 _33770_ (.A(_05583_),
    .B(_05585_),
    .X(_05587_));
 sky130_fd_sc_hd__or2_2 _33771_ (.A(_05586_),
    .B(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__a21oi_2 _33772_ (.A1(_05421_),
    .A2(_05425_),
    .B1(_05588_),
    .Y(_05589_));
 sky130_fd_sc_hd__and3_2 _33773_ (.A(_05588_),
    .B(_05421_),
    .C(_05425_),
    .X(_05591_));
 sky130_fd_sc_hd__nor2_2 _33774_ (.A(_05589_),
    .B(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__o21ai_2 _33775_ (.A1(_05404_),
    .A2(_05401_),
    .B1(_05400_),
    .Y(_05593_));
 sky130_fd_sc_hd__and2_2 _33776_ (.A(_05088_),
    .B(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__o21a_2 _33777_ (.A1(_05085_),
    .A2(_05403_),
    .B1(_05593_),
    .X(_05595_));
 sky130_fd_sc_hd__and2b_2 _33778_ (.A_N(_05396_),
    .B(_05393_),
    .X(_05596_));
 sky130_fd_sc_hd__and2b_2 _33779_ (.A_N(_05397_),
    .B(_05398_),
    .X(_05597_));
 sky130_fd_sc_hd__and2b_2 _33780_ (.A_N(_05391_),
    .B(_05392_),
    .X(_05598_));
 sky130_fd_sc_hd__inv_2 _33781_ (.A(_05386_),
    .Y(_05599_));
 sky130_fd_sc_hd__nand3_2 _33782_ (.A(_05008_),
    .B(_05289_),
    .C(_05290_),
    .Y(_05600_));
 sky130_fd_sc_hd__and4_2 _33783_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[59]),
    .D(iX[60]),
    .X(_05602_));
 sky130_fd_sc_hd__a22oi_2 _33784_ (.A1(iY[45]),
    .A2(iX[59]),
    .B1(iX[60]),
    .B2(iY[44]),
    .Y(_05603_));
 sky130_fd_sc_hd__nand2_2 _33785_ (.A(iY[46]),
    .B(iX[58]),
    .Y(_05604_));
 sky130_fd_sc_hd__o21a_2 _33786_ (.A1(_05602_),
    .A2(_05603_),
    .B1(_05604_),
    .X(_05605_));
 sky130_fd_sc_hd__nor3_2 _33787_ (.A(_05602_),
    .B(_05603_),
    .C(_05604_),
    .Y(_05606_));
 sky130_fd_sc_hd__nor2_2 _33788_ (.A(_05605_),
    .B(_05606_),
    .Y(_05607_));
 sky130_fd_sc_hd__inv_2 _33789_ (.A(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__and3_2 _33790_ (.A(iY[41]),
    .B(iX[61]),
    .C(_05274_),
    .X(_05609_));
 sky130_fd_sc_hd__and3_2 _33791_ (.A(iY[41]),
    .B(iX[63]),
    .C(_05274_),
    .X(_05610_));
 sky130_fd_sc_hd__a21o_2 _33792_ (.A1(iY[41]),
    .A2(iX[63]),
    .B1(_05274_),
    .X(_05611_));
 sky130_fd_sc_hd__and2b_2 _33793_ (.A_N(_05610_),
    .B(_05611_),
    .X(_05613_));
 sky130_fd_sc_hd__nand2_2 _33794_ (.A(iY[43]),
    .B(iX[61]),
    .Y(_05614_));
 sky130_fd_sc_hd__xnor2_2 _33795_ (.A(_05613_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__o21a_2 _33796_ (.A1(_05609_),
    .A2(_05279_),
    .B1(_05615_),
    .X(_05616_));
 sky130_fd_sc_hd__nor3_2 _33797_ (.A(_05609_),
    .B(_05279_),
    .C(_05615_),
    .Y(_05617_));
 sky130_fd_sc_hd__or2_2 _33798_ (.A(_05616_),
    .B(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__nor2_2 _33799_ (.A(_05608_),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__and2_2 _33800_ (.A(_05608_),
    .B(_05618_),
    .X(_05620_));
 sky130_fd_sc_hd__or2_2 _33801_ (.A(_05619_),
    .B(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__nor3_2 _33802_ (.A(_04239_),
    .B(_04980_),
    .C(_05621_),
    .Y(_05622_));
 sky130_fd_sc_hd__o21a_2 _33803_ (.A1(_04239_),
    .A2(_04980_),
    .B1(_05621_),
    .X(_05624_));
 sky130_fd_sc_hd__or2_2 _33804_ (.A(_05622_),
    .B(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__or3_2 _33805_ (.A(_05278_),
    .B(_05279_),
    .C(_05281_),
    .X(_05626_));
 sky130_fd_sc_hd__a21bo_2 _33806_ (.A1(_05272_),
    .A2(_05282_),
    .B1_N(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__xor2_2 _33807_ (.A(_05625_),
    .B(_05627_),
    .X(_05628_));
 sky130_fd_sc_hd__and2_2 _33808_ (.A(_05289_),
    .B(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__nor2_2 _33809_ (.A(_05289_),
    .B(_05628_),
    .Y(_05630_));
 sky130_fd_sc_hd__nor2_2 _33810_ (.A(_05629_),
    .B(_05630_),
    .Y(_05631_));
 sky130_fd_sc_hd__inv_2 _33811_ (.A(_05324_),
    .Y(_05632_));
 sky130_fd_sc_hd__or2b_2 _33812_ (.A(_05267_),
    .B_N(_05287_),
    .X(_05633_));
 sky130_fd_sc_hd__and4_2 _33813_ (.A(iX[50]),
    .B(iX[51]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_05635_));
 sky130_fd_sc_hd__a22oi_2 _33814_ (.A1(iX[51]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[50]),
    .Y(_05636_));
 sky130_fd_sc_hd__nor2_2 _33815_ (.A(_05635_),
    .B(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hd__nand2_2 _33816_ (.A(iX[49]),
    .B(iY[55]),
    .Y(_05638_));
 sky130_fd_sc_hd__xnor2_2 _33817_ (.A(_05637_),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__and4_2 _33818_ (.A(iY[50]),
    .B(iY[51]),
    .C(iX[53]),
    .D(iX[54]),
    .X(_05640_));
 sky130_fd_sc_hd__a22oi_2 _33819_ (.A1(iY[51]),
    .A2(iX[53]),
    .B1(iX[54]),
    .B2(iY[50]),
    .Y(_05641_));
 sky130_fd_sc_hd__nor2_2 _33820_ (.A(_05640_),
    .B(_05641_),
    .Y(_05642_));
 sky130_fd_sc_hd__nand2_2 _33821_ (.A(iX[52]),
    .B(iY[52]),
    .Y(_05643_));
 sky130_fd_sc_hd__xnor2_2 _33822_ (.A(_05642_),
    .B(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__o21ba_2 _33823_ (.A1(_05301_),
    .A2(_05303_),
    .B1_N(_05300_),
    .X(_05646_));
 sky130_fd_sc_hd__xnor2_2 _33824_ (.A(_05644_),
    .B(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__and2_2 _33825_ (.A(_05639_),
    .B(_05647_),
    .X(_05648_));
 sky130_fd_sc_hd__nor2_2 _33826_ (.A(_05639_),
    .B(_05647_),
    .Y(_05649_));
 sky130_fd_sc_hd__or2_2 _33827_ (.A(_05648_),
    .B(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__or3_2 _33828_ (.A(_05312_),
    .B(_05316_),
    .C(_05318_),
    .X(_05651_));
 sky130_fd_sc_hd__o21ba_2 _33829_ (.A1(_05269_),
    .A2(_05271_),
    .B1_N(_05268_),
    .X(_05652_));
 sky130_fd_sc_hd__and4_2 _33830_ (.A(iY[47]),
    .B(iY[48]),
    .C(iX[56]),
    .D(iX[57]),
    .X(_05653_));
 sky130_fd_sc_hd__a22oi_2 _33831_ (.A1(iY[48]),
    .A2(iX[56]),
    .B1(iX[57]),
    .B2(iY[47]),
    .Y(_05654_));
 sky130_fd_sc_hd__nor2_2 _33832_ (.A(_05653_),
    .B(_05654_),
    .Y(_05655_));
 sky130_fd_sc_hd__nand2_2 _33833_ (.A(iY[49]),
    .B(iX[55]),
    .Y(_05657_));
 sky130_fd_sc_hd__xnor2_2 _33834_ (.A(_05655_),
    .B(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__xnor2_2 _33835_ (.A(_05652_),
    .B(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__o21ai_2 _33836_ (.A1(_05313_),
    .A2(_05318_),
    .B1(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__or3_2 _33837_ (.A(_05313_),
    .B(_05318_),
    .C(_05659_),
    .X(_05661_));
 sky130_fd_sc_hd__nand2_2 _33838_ (.A(_05660_),
    .B(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hd__a21oi_2 _33839_ (.A1(_05651_),
    .A2(_05321_),
    .B1(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__and3_2 _33840_ (.A(_05651_),
    .B(_05321_),
    .C(_05662_),
    .X(_05664_));
 sky130_fd_sc_hd__or3_2 _33841_ (.A(_05650_),
    .B(_05663_),
    .C(_05664_),
    .X(_05665_));
 sky130_fd_sc_hd__o21ai_2 _33842_ (.A1(_05663_),
    .A2(_05664_),
    .B1(_05650_),
    .Y(_05666_));
 sky130_fd_sc_hd__nand2_2 _33843_ (.A(_05665_),
    .B(_05666_),
    .Y(_05668_));
 sky130_fd_sc_hd__a21oi_2 _33844_ (.A1(_05285_),
    .A2(_05633_),
    .B1(_05668_),
    .Y(_05669_));
 sky130_fd_sc_hd__and3_2 _33845_ (.A(_05285_),
    .B(_05633_),
    .C(_05668_),
    .X(_05670_));
 sky130_fd_sc_hd__a211o_2 _33846_ (.A1(_05632_),
    .A2(_05326_),
    .B1(_05669_),
    .C1(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__o211ai_2 _33847_ (.A1(_05669_),
    .A2(_05670_),
    .B1(_05632_),
    .C1(_05326_),
    .Y(_05672_));
 sky130_fd_sc_hd__and3_2 _33848_ (.A(_05631_),
    .B(_05671_),
    .C(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__a21oi_2 _33849_ (.A1(_05671_),
    .A2(_05672_),
    .B1(_05631_),
    .Y(_05674_));
 sky130_fd_sc_hd__a211o_2 _33850_ (.A1(_05600_),
    .A2(_05334_),
    .B1(_05673_),
    .C1(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__o211ai_2 _33851_ (.A1(_05673_),
    .A2(_05674_),
    .B1(_05600_),
    .C1(_05334_),
    .Y(_05676_));
 sky130_fd_sc_hd__inv_2 _33852_ (.A(_05378_),
    .Y(_05677_));
 sky130_fd_sc_hd__or2b_2 _33853_ (.A(_05330_),
    .B_N(_05332_),
    .X(_05679_));
 sky130_fd_sc_hd__inv_2 _33854_ (.A(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__and4_2 _33855_ (.A(iX[44]),
    .B(iX[45]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_05681_));
 sky130_fd_sc_hd__a22oi_2 _33856_ (.A1(iX[45]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[44]),
    .Y(_05682_));
 sky130_fd_sc_hd__nor2_2 _33857_ (.A(_05681_),
    .B(_05682_),
    .Y(_05683_));
 sky130_fd_sc_hd__nand2_2 _33858_ (.A(iX[43]),
    .B(iY[61]),
    .Y(_05684_));
 sky130_fd_sc_hd__xnor2_2 _33859_ (.A(_05683_),
    .B(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__o21ba_2 _33860_ (.A1(_05343_),
    .A2(_05345_),
    .B1_N(_05342_),
    .X(_05686_));
 sky130_fd_sc_hd__xnor2_2 _33861_ (.A(_05685_),
    .B(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__and2_2 _33862_ (.A(iX[42]),
    .B(iY[62]),
    .X(_05688_));
 sky130_fd_sc_hd__or2_2 _33863_ (.A(_05687_),
    .B(_05688_),
    .X(_05690_));
 sky130_fd_sc_hd__nand2_2 _33864_ (.A(_05687_),
    .B(_05688_),
    .Y(_05691_));
 sky130_fd_sc_hd__and2b_2 _33865_ (.A_N(_05347_),
    .B(_05346_),
    .X(_05692_));
 sky130_fd_sc_hd__a31o_2 _33866_ (.A1(iX[41]),
    .A2(iY[62]),
    .A3(_05348_),
    .B1(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__nand3_2 _33867_ (.A(_05690_),
    .B(_05691_),
    .C(_05693_),
    .Y(_05694_));
 sky130_fd_sc_hd__a21o_2 _33868_ (.A1(_05690_),
    .A2(_05691_),
    .B1(_05693_),
    .X(_05695_));
 sky130_fd_sc_hd__nand2_2 _33869_ (.A(_05694_),
    .B(_05695_),
    .Y(_05696_));
 sky130_fd_sc_hd__nand2_2 _33870_ (.A(iX[41]),
    .B(iY[63]),
    .Y(_05697_));
 sky130_fd_sc_hd__nand2_2 _33871_ (.A(_05696_),
    .B(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__or2_2 _33872_ (.A(_05696_),
    .B(_05697_),
    .X(_05699_));
 sky130_fd_sc_hd__and2_2 _33873_ (.A(_05698_),
    .B(_05699_),
    .X(_05701_));
 sky130_fd_sc_hd__or2b_2 _33874_ (.A(_05362_),
    .B_N(_05367_),
    .X(_05702_));
 sky130_fd_sc_hd__or2b_2 _33875_ (.A(_05360_),
    .B_N(_05368_),
    .X(_05703_));
 sky130_fd_sc_hd__and2b_2 _33876_ (.A_N(_05305_),
    .B(_05304_),
    .X(_05704_));
 sky130_fd_sc_hd__o21ba_2 _33877_ (.A1(_05364_),
    .A2(_05366_),
    .B1_N(_05363_),
    .X(_05705_));
 sky130_fd_sc_hd__o21ba_2 _33878_ (.A1(_05296_),
    .A2(_05298_),
    .B1_N(_05294_),
    .X(_05706_));
 sky130_fd_sc_hd__and4_2 _33879_ (.A(iX[47]),
    .B(iX[48]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_05707_));
 sky130_fd_sc_hd__a22oi_2 _33880_ (.A1(iX[48]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[47]),
    .Y(_05708_));
 sky130_fd_sc_hd__nor2_2 _33881_ (.A(_05707_),
    .B(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__nand2_2 _33882_ (.A(iX[46]),
    .B(iY[58]),
    .Y(_05710_));
 sky130_fd_sc_hd__xnor2_2 _33883_ (.A(_05709_),
    .B(_05710_),
    .Y(_05712_));
 sky130_fd_sc_hd__xnor2_2 _33884_ (.A(_05706_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__xnor2_2 _33885_ (.A(_05705_),
    .B(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__o21a_2 _33886_ (.A1(_05704_),
    .A2(_05308_),
    .B1(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__nor3_2 _33887_ (.A(_05704_),
    .B(_05308_),
    .C(_05714_),
    .Y(_05716_));
 sky130_fd_sc_hd__a211oi_2 _33888_ (.A1(_05702_),
    .A2(_05703_),
    .B1(_05715_),
    .C1(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__o211a_2 _33889_ (.A1(_05715_),
    .A2(_05716_),
    .B1(_05702_),
    .C1(_05703_),
    .X(_05718_));
 sky130_fd_sc_hd__nor2_2 _33890_ (.A(_05370_),
    .B(_05373_),
    .Y(_05719_));
 sky130_fd_sc_hd__or3_2 _33891_ (.A(_05717_),
    .B(_05718_),
    .C(_05719_),
    .X(_05720_));
 sky130_fd_sc_hd__o21ai_2 _33892_ (.A1(_05717_),
    .A2(_05718_),
    .B1(_05719_),
    .Y(_05721_));
 sky130_fd_sc_hd__and3_2 _33893_ (.A(_05701_),
    .B(_05720_),
    .C(_05721_),
    .X(_05723_));
 sky130_fd_sc_hd__a21oi_2 _33894_ (.A1(_05720_),
    .A2(_05721_),
    .B1(_05701_),
    .Y(_05724_));
 sky130_fd_sc_hd__or3_2 _33895_ (.A(_05680_),
    .B(_05723_),
    .C(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__o21ai_2 _33896_ (.A1(_05723_),
    .A2(_05724_),
    .B1(_05680_),
    .Y(_05726_));
 sky130_fd_sc_hd__nand2_2 _33897_ (.A(_05725_),
    .B(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__a21o_2 _33898_ (.A1(_05376_),
    .A2(_05677_),
    .B1(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__nand3_2 _33899_ (.A(_05376_),
    .B(_05677_),
    .C(_05727_),
    .Y(_05729_));
 sky130_fd_sc_hd__nand4_2 _33900_ (.A(_05675_),
    .B(_05676_),
    .C(_05728_),
    .D(_05729_),
    .Y(_05730_));
 sky130_fd_sc_hd__a22o_2 _33901_ (.A1(_05675_),
    .A2(_05676_),
    .B1(_05728_),
    .B2(_05729_),
    .X(_05731_));
 sky130_fd_sc_hd__o211a_2 _33902_ (.A1(_05337_),
    .A2(_05599_),
    .B1(_05730_),
    .C1(_05731_),
    .X(_05732_));
 sky130_fd_sc_hd__a211oi_2 _33903_ (.A1(_05730_),
    .A2(_05731_),
    .B1(_05337_),
    .C1(_05599_),
    .Y(_05734_));
 sky130_fd_sc_hd__or2_2 _33904_ (.A(_05732_),
    .B(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__nand2_2 _33905_ (.A(_05381_),
    .B(_05384_),
    .Y(_05736_));
 sky130_fd_sc_hd__xnor2_2 _33906_ (.A(_05735_),
    .B(_05736_),
    .Y(_05737_));
 sky130_fd_sc_hd__o21a_2 _33907_ (.A1(_05389_),
    .A2(_05598_),
    .B1(_05737_),
    .X(_05738_));
 sky130_fd_sc_hd__nor3_2 _33908_ (.A(_05389_),
    .B(_05598_),
    .C(_05737_),
    .Y(_05739_));
 sky130_fd_sc_hd__nor2_2 _33909_ (.A(_05738_),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__a31o_2 _33910_ (.A1(iX[40]),
    .A2(iY[63]),
    .A3(_05354_),
    .B1(_05352_),
    .X(_05741_));
 sky130_fd_sc_hd__xnor2_2 _33911_ (.A(_05740_),
    .B(_05741_),
    .Y(_05742_));
 sky130_fd_sc_hd__o21bai_2 _33912_ (.A1(_05596_),
    .A2(_05597_),
    .B1_N(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__or3b_2 _33913_ (.A(_05596_),
    .B(_05597_),
    .C_N(_05742_),
    .X(_05745_));
 sky130_fd_sc_hd__nand2_2 _33914_ (.A(_05743_),
    .B(_05745_),
    .Y(_05746_));
 sky130_fd_sc_hd__a211o_2 _33915_ (.A1(_05086_),
    .A2(_05594_),
    .B1(_05595_),
    .C1(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__a21o_2 _33916_ (.A1(_05086_),
    .A2(_05594_),
    .B1(_05595_),
    .X(_05748_));
 sky130_fd_sc_hd__nand2_2 _33917_ (.A(_05746_),
    .B(_05748_),
    .Y(_05749_));
 sky130_fd_sc_hd__and2_2 _33918_ (.A(_05747_),
    .B(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__buf_1 _33919_ (.A(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__xnor2_2 _33920_ (.A(_05592_),
    .B(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__nand2_2 _33921_ (.A(_13229_),
    .B(_05752_),
    .Y(_05753_));
 sky130_fd_sc_hd__or2_2 _33922_ (.A(_13229_),
    .B(_05752_),
    .X(_05754_));
 sky130_fd_sc_hd__nand2_2 _33923_ (.A(_05753_),
    .B(_05754_),
    .Y(_05756_));
 sky130_fd_sc_hd__and2_2 _33924_ (.A(_05409_),
    .B(_05410_),
    .X(_05757_));
 sky130_fd_sc_hd__xor2_2 _33925_ (.A(_05756_),
    .B(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__nor2_2 _33926_ (.A(_04759_),
    .B(_04760_),
    .Y(_05759_));
 sky130_fd_sc_hd__and3_2 _33927_ (.A(_05095_),
    .B(_05414_),
    .C(_05415_),
    .X(_05760_));
 sky130_fd_sc_hd__and4b_2 _33928_ (.A_N(_04415_),
    .B(_04416_),
    .C(_05759_),
    .D(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__and4b_2 _33929_ (.A_N(_04415_),
    .B(_04421_),
    .C(_05759_),
    .D(_05760_),
    .X(_05762_));
 sky130_fd_sc_hd__o21ba_2 _33930_ (.A1(_04413_),
    .A2(_04759_),
    .B1_N(_04760_),
    .X(_05763_));
 sky130_fd_sc_hd__a21bo_2 _33931_ (.A1(_05106_),
    .A2(_05414_),
    .B1_N(_05415_),
    .X(_05764_));
 sky130_fd_sc_hd__a21o_2 _33932_ (.A1(_05763_),
    .A2(_05760_),
    .B1(_05764_),
    .X(_05765_));
 sky130_fd_sc_hd__a211oi_2 _33933_ (.A1(_03682_),
    .A2(_05761_),
    .B1(_05762_),
    .C1(_05765_),
    .Y(_05767_));
 sky130_fd_sc_hd__xnor2_2 _33934_ (.A(_05758_),
    .B(_05767_),
    .Y(_05768_));
 sky130_fd_sc_hd__and2_2 _33935_ (.A(_13341_),
    .B(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__nor2_2 _33936_ (.A(_13341_),
    .B(_05768_),
    .Y(_05770_));
 sky130_fd_sc_hd__nor2_2 _33937_ (.A(_05769_),
    .B(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__or2_2 _33938_ (.A(_05102_),
    .B(_05419_),
    .X(_05772_));
 sky130_fd_sc_hd__or4b_2 _33939_ (.A(_04426_),
    .B(_05772_),
    .C(_04765_),
    .D_N(_05103_),
    .X(_05773_));
 sky130_fd_sc_hd__nor2_2 _33940_ (.A(_04427_),
    .B(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__inv_2 _33941_ (.A(_05104_),
    .Y(_05775_));
 sky130_fd_sc_hd__or2b_2 _33942_ (.A(_05418_),
    .B_N(_12911_),
    .X(_05776_));
 sky130_fd_sc_hd__and2b_2 _33943_ (.A_N(_12911_),
    .B(_05418_),
    .X(_05778_));
 sky130_fd_sc_hd__a21o_2 _33944_ (.A1(_05100_),
    .A2(_05776_),
    .B1(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__o221ai_2 _33945_ (.A1(_05775_),
    .A2(_05772_),
    .B1(_05773_),
    .B2(_04430_),
    .C1(_05779_),
    .Y(_05780_));
 sky130_fd_sc_hd__a21o_2 _33946_ (.A1(_03690_),
    .A2(_05774_),
    .B1(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__a21oi_2 _33947_ (.A1(_03689_),
    .A2(_05774_),
    .B1(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__xnor2_2 _33948_ (.A(_05771_),
    .B(_05782_),
    .Y(oO[72]));
 sky130_fd_sc_hd__and2b_2 _33949_ (.A_N(_05735_),
    .B(_05736_),
    .X(_05783_));
 sky130_fd_sc_hd__and3_2 _33950_ (.A(iY[43]),
    .B(iX[63]),
    .C(_05274_),
    .X(_05784_));
 sky130_fd_sc_hd__a22oi_2 _33951_ (.A1(iY[43]),
    .A2(iX[62]),
    .B1(iX[63]),
    .B2(iY[42]),
    .Y(_05785_));
 sky130_fd_sc_hd__or2_2 _33952_ (.A(_05784_),
    .B(_05785_),
    .X(_05786_));
 sky130_fd_sc_hd__a31o_2 _33953_ (.A1(iY[43]),
    .A2(iX[61]),
    .A3(_05611_),
    .B1(_05610_),
    .X(_05788_));
 sky130_fd_sc_hd__xnor2_2 _33954_ (.A(_05786_),
    .B(_05788_),
    .Y(_05789_));
 sky130_fd_sc_hd__and4_2 _33955_ (.A(iY[44]),
    .B(iY[45]),
    .C(iX[60]),
    .D(iX[61]),
    .X(_05790_));
 sky130_fd_sc_hd__a22oi_2 _33956_ (.A1(iY[45]),
    .A2(iX[60]),
    .B1(iX[61]),
    .B2(iY[44]),
    .Y(_05791_));
 sky130_fd_sc_hd__nor2_2 _33957_ (.A(_05790_),
    .B(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__nand2_2 _33958_ (.A(iY[46]),
    .B(iX[59]),
    .Y(_05793_));
 sky130_fd_sc_hd__xnor2_2 _33959_ (.A(_05792_),
    .B(_05793_),
    .Y(_05794_));
 sky130_fd_sc_hd__xor2_2 _33960_ (.A(_05789_),
    .B(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__o21a_2 _33961_ (.A1(_05616_),
    .A2(_05619_),
    .B1(_05795_),
    .X(_05796_));
 sky130_fd_sc_hd__nor3_2 _33962_ (.A(_05616_),
    .B(_05619_),
    .C(_05795_),
    .Y(_05797_));
 sky130_fd_sc_hd__or2_2 _33963_ (.A(_05796_),
    .B(_05797_),
    .X(_05799_));
 sky130_fd_sc_hd__inv_2 _33964_ (.A(_05663_),
    .Y(_05800_));
 sky130_fd_sc_hd__and2b_2 _33965_ (.A_N(_05625_),
    .B(_05627_),
    .X(_05801_));
 sky130_fd_sc_hd__and4_2 _33966_ (.A(iX[51]),
    .B(iX[52]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_05802_));
 sky130_fd_sc_hd__a22oi_2 _33967_ (.A1(iX[52]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[51]),
    .Y(_05803_));
 sky130_fd_sc_hd__nor2_2 _33968_ (.A(_05802_),
    .B(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__nand2_2 _33969_ (.A(iX[50]),
    .B(iY[55]),
    .Y(_05805_));
 sky130_fd_sc_hd__xnor2_2 _33970_ (.A(_05804_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__and4_2 _33971_ (.A(iY[50]),
    .B(iY[51]),
    .C(iX[54]),
    .D(iX[55]),
    .X(_05807_));
 sky130_fd_sc_hd__a22oi_2 _33972_ (.A1(iY[51]),
    .A2(iX[54]),
    .B1(iX[55]),
    .B2(iY[50]),
    .Y(_05808_));
 sky130_fd_sc_hd__nor2_2 _33973_ (.A(_05807_),
    .B(_05808_),
    .Y(_05810_));
 sky130_fd_sc_hd__nand2_2 _33974_ (.A(iY[52]),
    .B(iX[53]),
    .Y(_05811_));
 sky130_fd_sc_hd__xnor2_2 _33975_ (.A(_05810_),
    .B(_05811_),
    .Y(_05812_));
 sky130_fd_sc_hd__o21ba_2 _33976_ (.A1(_05641_),
    .A2(_05643_),
    .B1_N(_05640_),
    .X(_05813_));
 sky130_fd_sc_hd__xnor2_2 _33977_ (.A(_05812_),
    .B(_05813_),
    .Y(_05814_));
 sky130_fd_sc_hd__and2_2 _33978_ (.A(_05806_),
    .B(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__nor2_2 _33979_ (.A(_05806_),
    .B(_05814_),
    .Y(_05816_));
 sky130_fd_sc_hd__or2_2 _33980_ (.A(_05815_),
    .B(_05816_),
    .X(_05817_));
 sky130_fd_sc_hd__or2b_2 _33981_ (.A(_05652_),
    .B_N(_05658_),
    .X(_05818_));
 sky130_fd_sc_hd__a31o_2 _33982_ (.A1(iY[49]),
    .A2(iX[55]),
    .A3(_05655_),
    .B1(_05653_),
    .X(_05819_));
 sky130_fd_sc_hd__and4_2 _33983_ (.A(iY[47]),
    .B(iY[48]),
    .C(iX[57]),
    .D(iX[58]),
    .X(_05821_));
 sky130_fd_sc_hd__a22oi_2 _33984_ (.A1(iY[48]),
    .A2(iX[57]),
    .B1(iX[58]),
    .B2(iY[47]),
    .Y(_05822_));
 sky130_fd_sc_hd__nand2_2 _33985_ (.A(iY[49]),
    .B(iX[56]),
    .Y(_05823_));
 sky130_fd_sc_hd__o21a_2 _33986_ (.A1(_05821_),
    .A2(_05822_),
    .B1(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__nor3_2 _33987_ (.A(_05821_),
    .B(_05822_),
    .C(_05823_),
    .Y(_05825_));
 sky130_fd_sc_hd__nor2_2 _33988_ (.A(_05824_),
    .B(_05825_),
    .Y(_05826_));
 sky130_fd_sc_hd__o21ai_2 _33989_ (.A1(_05602_),
    .A2(_05606_),
    .B1(_05826_),
    .Y(_05827_));
 sky130_fd_sc_hd__or3_2 _33990_ (.A(_05602_),
    .B(_05606_),
    .C(_05826_),
    .X(_05828_));
 sky130_fd_sc_hd__and2_2 _33991_ (.A(_05827_),
    .B(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__xnor2_2 _33992_ (.A(_05819_),
    .B(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__a21oi_2 _33993_ (.A1(_05818_),
    .A2(_05660_),
    .B1(_05830_),
    .Y(_05832_));
 sky130_fd_sc_hd__and3_2 _33994_ (.A(_05818_),
    .B(_05660_),
    .C(_05830_),
    .X(_05833_));
 sky130_fd_sc_hd__or3_2 _33995_ (.A(_05817_),
    .B(_05832_),
    .C(_05833_),
    .X(_05834_));
 sky130_fd_sc_hd__o21ai_2 _33996_ (.A1(_05832_),
    .A2(_05833_),
    .B1(_05817_),
    .Y(_05835_));
 sky130_fd_sc_hd__o211a_2 _33997_ (.A1(_05622_),
    .A2(_05801_),
    .B1(_05834_),
    .C1(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__a211oi_2 _33998_ (.A1(_05834_),
    .A2(_05835_),
    .B1(_05622_),
    .C1(_05801_),
    .Y(_05837_));
 sky130_fd_sc_hd__a211oi_2 _33999_ (.A1(_05800_),
    .A2(_05665_),
    .B1(_05836_),
    .C1(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__o211a_2 _34000_ (.A1(_05836_),
    .A2(_05837_),
    .B1(_05800_),
    .C1(_05665_),
    .X(_05839_));
 sky130_fd_sc_hd__or3_2 _34001_ (.A(_05799_),
    .B(_05838_),
    .C(_05839_),
    .X(_05840_));
 sky130_fd_sc_hd__o21ai_2 _34002_ (.A1(_05838_),
    .A2(_05839_),
    .B1(_05799_),
    .Y(_05841_));
 sky130_fd_sc_hd__o211ai_2 _34003_ (.A1(_05630_),
    .A2(_05673_),
    .B1(_05840_),
    .C1(_05841_),
    .Y(_05843_));
 sky130_fd_sc_hd__a211o_2 _34004_ (.A1(_05840_),
    .A2(_05841_),
    .B1(_05630_),
    .C1(_05673_),
    .X(_05844_));
 sky130_fd_sc_hd__inv_2 _34005_ (.A(_05723_),
    .Y(_05845_));
 sky130_fd_sc_hd__or2b_2 _34006_ (.A(_05669_),
    .B_N(_05671_),
    .X(_05846_));
 sky130_fd_sc_hd__inv_2 _34007_ (.A(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__or2b_2 _34008_ (.A(_05686_),
    .B_N(_05685_),
    .X(_05848_));
 sky130_fd_sc_hd__and4_2 _34009_ (.A(iX[45]),
    .B(iX[46]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_05849_));
 sky130_fd_sc_hd__a22oi_2 _34010_ (.A1(iX[46]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[45]),
    .Y(_05850_));
 sky130_fd_sc_hd__nor2_2 _34011_ (.A(_05849_),
    .B(_05850_),
    .Y(_05851_));
 sky130_fd_sc_hd__nand2_2 _34012_ (.A(iX[44]),
    .B(iY[61]),
    .Y(_05852_));
 sky130_fd_sc_hd__xnor2_2 _34013_ (.A(_05851_),
    .B(_05852_),
    .Y(_05854_));
 sky130_fd_sc_hd__o21ba_2 _34014_ (.A1(_05682_),
    .A2(_05684_),
    .B1_N(_05681_),
    .X(_05855_));
 sky130_fd_sc_hd__xnor2_2 _34015_ (.A(_05854_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__nand2_2 _34016_ (.A(iX[43]),
    .B(iY[62]),
    .Y(_05857_));
 sky130_fd_sc_hd__xor2_2 _34017_ (.A(_05856_),
    .B(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__a21oi_2 _34018_ (.A1(_05848_),
    .A2(_05691_),
    .B1(_05858_),
    .Y(_05859_));
 sky130_fd_sc_hd__and3_2 _34019_ (.A(_05848_),
    .B(_05691_),
    .C(_05858_),
    .X(_05860_));
 sky130_fd_sc_hd__nor2_2 _34020_ (.A(_05859_),
    .B(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__a21oi_2 _34021_ (.A1(iX[42]),
    .A2(iY[63]),
    .B1(_05861_),
    .Y(_05862_));
 sky130_fd_sc_hd__and3_2 _34022_ (.A(iX[42]),
    .B(iY[63]),
    .C(_05861_),
    .X(_05863_));
 sky130_fd_sc_hd__nor2_2 _34023_ (.A(_05862_),
    .B(_05863_),
    .Y(_05865_));
 sky130_fd_sc_hd__or2b_2 _34024_ (.A(_05706_),
    .B_N(_05712_),
    .X(_05866_));
 sky130_fd_sc_hd__or2b_2 _34025_ (.A(_05705_),
    .B_N(_05713_),
    .X(_05867_));
 sky130_fd_sc_hd__and2b_2 _34026_ (.A_N(_05646_),
    .B(_05644_),
    .X(_05868_));
 sky130_fd_sc_hd__o21ba_2 _34027_ (.A1(_05708_),
    .A2(_05710_),
    .B1_N(_05707_),
    .X(_05869_));
 sky130_fd_sc_hd__o21ba_2 _34028_ (.A1(_05636_),
    .A2(_05638_),
    .B1_N(_05635_),
    .X(_05870_));
 sky130_fd_sc_hd__and4_2 _34029_ (.A(iX[48]),
    .B(iX[49]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_05871_));
 sky130_fd_sc_hd__a22oi_2 _34030_ (.A1(iX[49]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[48]),
    .Y(_05872_));
 sky130_fd_sc_hd__nor2_2 _34031_ (.A(_05871_),
    .B(_05872_),
    .Y(_05873_));
 sky130_fd_sc_hd__nand2_2 _34032_ (.A(iX[47]),
    .B(iY[58]),
    .Y(_05874_));
 sky130_fd_sc_hd__xnor2_2 _34033_ (.A(_05873_),
    .B(_05874_),
    .Y(_05876_));
 sky130_fd_sc_hd__xnor2_2 _34034_ (.A(_05870_),
    .B(_05876_),
    .Y(_05877_));
 sky130_fd_sc_hd__xnor2_2 _34035_ (.A(_05869_),
    .B(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__o21a_2 _34036_ (.A1(_05868_),
    .A2(_05648_),
    .B1(_05878_),
    .X(_05879_));
 sky130_fd_sc_hd__nor3_2 _34037_ (.A(_05868_),
    .B(_05648_),
    .C(_05878_),
    .Y(_05880_));
 sky130_fd_sc_hd__a211oi_2 _34038_ (.A1(_05866_),
    .A2(_05867_),
    .B1(_05879_),
    .C1(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__o211a_2 _34039_ (.A1(_05879_),
    .A2(_05880_),
    .B1(_05866_),
    .C1(_05867_),
    .X(_05882_));
 sky130_fd_sc_hd__nor2_2 _34040_ (.A(_05715_),
    .B(_05717_),
    .Y(_05883_));
 sky130_fd_sc_hd__or3_2 _34041_ (.A(_05881_),
    .B(_05882_),
    .C(_05883_),
    .X(_05884_));
 sky130_fd_sc_hd__o21ai_2 _34042_ (.A1(_05881_),
    .A2(_05882_),
    .B1(_05883_),
    .Y(_05885_));
 sky130_fd_sc_hd__and3_2 _34043_ (.A(_05865_),
    .B(_05884_),
    .C(_05885_),
    .X(_05887_));
 sky130_fd_sc_hd__a21oi_2 _34044_ (.A1(_05884_),
    .A2(_05885_),
    .B1(_05865_),
    .Y(_05888_));
 sky130_fd_sc_hd__or3_2 _34045_ (.A(_05847_),
    .B(_05887_),
    .C(_05888_),
    .X(_05889_));
 sky130_fd_sc_hd__o21ai_2 _34046_ (.A1(_05887_),
    .A2(_05888_),
    .B1(_05847_),
    .Y(_05890_));
 sky130_fd_sc_hd__nand2_2 _34047_ (.A(_05889_),
    .B(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__a21o_2 _34048_ (.A1(_05720_),
    .A2(_05845_),
    .B1(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__nand3_2 _34049_ (.A(_05720_),
    .B(_05845_),
    .C(_05891_),
    .Y(_05893_));
 sky130_fd_sc_hd__nand4_2 _34050_ (.A(_05843_),
    .B(_05844_),
    .C(_05892_),
    .D(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__a22o_2 _34051_ (.A1(_05843_),
    .A2(_05844_),
    .B1(_05892_),
    .B2(_05893_),
    .X(_05895_));
 sky130_fd_sc_hd__nand2_2 _34052_ (.A(_05675_),
    .B(_05730_),
    .Y(_05896_));
 sky130_fd_sc_hd__and3_2 _34053_ (.A(_05894_),
    .B(_05895_),
    .C(_05896_),
    .X(_05898_));
 sky130_fd_sc_hd__a21oi_2 _34054_ (.A1(_05894_),
    .A2(_05895_),
    .B1(_05896_),
    .Y(_05899_));
 sky130_fd_sc_hd__a211oi_2 _34055_ (.A1(_05725_),
    .A2(_05728_),
    .B1(_05898_),
    .C1(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__o211a_2 _34056_ (.A1(_05898_),
    .A2(_05899_),
    .B1(_05725_),
    .C1(_05728_),
    .X(_05901_));
 sky130_fd_sc_hd__nor2_2 _34057_ (.A(_05900_),
    .B(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__o21a_2 _34058_ (.A1(_05732_),
    .A2(_05783_),
    .B1(_05902_),
    .X(_05903_));
 sky130_fd_sc_hd__nor3_2 _34059_ (.A(_05732_),
    .B(_05783_),
    .C(_05902_),
    .Y(_05904_));
 sky130_fd_sc_hd__a211oi_2 _34060_ (.A1(_05694_),
    .A2(_05699_),
    .B1(_05903_),
    .C1(_05904_),
    .Y(_05905_));
 sky130_fd_sc_hd__o211a_2 _34061_ (.A1(_05903_),
    .A2(_05904_),
    .B1(_05694_),
    .C1(_05699_),
    .X(_05906_));
 sky130_fd_sc_hd__nor2_2 _34062_ (.A(_05905_),
    .B(_05906_),
    .Y(_05907_));
 sky130_fd_sc_hd__a21o_2 _34063_ (.A1(_05740_),
    .A2(_05741_),
    .B1(_05738_),
    .X(_05909_));
 sky130_fd_sc_hd__xnor2_2 _34064_ (.A(_05907_),
    .B(_05909_),
    .Y(_05910_));
 sky130_fd_sc_hd__and2_2 _34065_ (.A(_05743_),
    .B(_05747_),
    .X(_05911_));
 sky130_fd_sc_hd__xor2_2 _34066_ (.A(_05910_),
    .B(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__o21a_2 _34067_ (.A1(_05430_),
    .A2(_05431_),
    .B1(_05429_),
    .X(_05913_));
 sky130_fd_sc_hd__or2b_2 _34068_ (.A(_05488_),
    .B_N(_05439_),
    .X(_05914_));
 sky130_fd_sc_hd__or2b_2 _34069_ (.A(_05489_),
    .B_N(_05436_),
    .X(_05915_));
 sky130_fd_sc_hd__and2b_2 _34070_ (.A_N(_05462_),
    .B(_05463_),
    .X(_05916_));
 sky130_fd_sc_hd__and2b_2 _34071_ (.A_N(_05443_),
    .B(_05464_),
    .X(_05917_));
 sky130_fd_sc_hd__nor2_2 _34072_ (.A(_05916_),
    .B(_05917_),
    .Y(_05918_));
 sky130_fd_sc_hd__a21oi_2 _34073_ (.A1(_05914_),
    .A2(_05915_),
    .B1(_05918_),
    .Y(_05920_));
 sky130_fd_sc_hd__and3_2 _34074_ (.A(_05914_),
    .B(_05915_),
    .C(_05918_),
    .X(_05921_));
 sky130_fd_sc_hd__nor2_2 _34075_ (.A(_05920_),
    .B(_05921_),
    .Y(_05922_));
 sky130_fd_sc_hd__a21o_2 _34076_ (.A1(_05465_),
    .A2(_05487_),
    .B1(_05485_),
    .X(_05923_));
 sky130_fd_sc_hd__or2b_2 _34077_ (.A(_05530_),
    .B_N(_05494_),
    .X(_05924_));
 sky130_fd_sc_hd__or2b_2 _34078_ (.A(_05491_),
    .B_N(_05531_),
    .X(_05925_));
 sky130_fd_sc_hd__nand2_2 _34079_ (.A(_05924_),
    .B(_05925_),
    .Y(_05926_));
 sky130_fd_sc_hd__o31a_2 _34080_ (.A1(_16288_),
    .A2(_05440_),
    .A3(_05446_),
    .B1(_05444_),
    .X(_05927_));
 sky130_fd_sc_hd__nand2_2 _34081_ (.A(_15888_),
    .B(_01522_),
    .Y(_05928_));
 sky130_fd_sc_hd__or3_2 _34082_ (.A(_01576_),
    .B(_02317_),
    .C(_05928_),
    .X(_05929_));
 sky130_fd_sc_hd__buf_1 _34083_ (.A(_02317_),
    .X(_05931_));
 sky130_fd_sc_hd__o21ai_2 _34084_ (.A1(_01576_),
    .A2(_05931_),
    .B1(_05928_),
    .Y(_05932_));
 sky130_fd_sc_hd__nand2_2 _34085_ (.A(_05929_),
    .B(_05932_),
    .Y(_05933_));
 sky130_fd_sc_hd__nor2_2 _34086_ (.A(_01797_),
    .B(_03318_),
    .Y(_05934_));
 sky130_fd_sc_hd__xnor2_2 _34087_ (.A(_05933_),
    .B(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__nand2_2 _34088_ (.A(_02989_),
    .B(_01757_),
    .Y(_05936_));
 sky130_fd_sc_hd__xnor2_2 _34089_ (.A(_05452_),
    .B(_05936_),
    .Y(_05937_));
 sky130_fd_sc_hd__nand2_2 _34090_ (.A(_02983_),
    .B(_03327_),
    .Y(_05938_));
 sky130_fd_sc_hd__xnor2_2 _34091_ (.A(_05937_),
    .B(_05938_),
    .Y(_05939_));
 sky130_fd_sc_hd__o22a_2 _34092_ (.A1(_05451_),
    .A2(_05452_),
    .B1(_05454_),
    .B2(_05455_),
    .X(_05940_));
 sky130_fd_sc_hd__nor2_2 _34093_ (.A(_05939_),
    .B(_05940_),
    .Y(_05942_));
 sky130_fd_sc_hd__and2_2 _34094_ (.A(_05939_),
    .B(_05940_),
    .X(_05943_));
 sky130_fd_sc_hd__nor2_2 _34095_ (.A(_05942_),
    .B(_05943_),
    .Y(_05944_));
 sky130_fd_sc_hd__xnor2_2 _34096_ (.A(_05935_),
    .B(_05944_),
    .Y(_05945_));
 sky130_fd_sc_hd__a21o_2 _34097_ (.A1(_05449_),
    .A2(_05460_),
    .B1(_05458_),
    .X(_05946_));
 sky130_fd_sc_hd__xnor2_2 _34098_ (.A(_05945_),
    .B(_05946_),
    .Y(_05947_));
 sky130_fd_sc_hd__xnor2_2 _34099_ (.A(_05927_),
    .B(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__and2b_2 _34100_ (.A_N(_05479_),
    .B(_05474_),
    .X(_05949_));
 sky130_fd_sc_hd__a21oi_2 _34101_ (.A1(_05473_),
    .A2(_05480_),
    .B1(_05949_),
    .Y(_05950_));
 sky130_fd_sc_hd__o21a_2 _34102_ (.A1(_05502_),
    .A2(_05513_),
    .B1(_05511_),
    .X(_05951_));
 sky130_fd_sc_hd__a2bb2o_2 _34103_ (.A1_N(_05475_),
    .A2_N(_05476_),
    .B1(_05477_),
    .B2(_05478_),
    .X(_05953_));
 sky130_fd_sc_hd__nand2_2 _34104_ (.A(_05496_),
    .B(_05501_),
    .Y(_05954_));
 sky130_fd_sc_hd__nor3_2 _34105_ (.A(_04504_),
    .B(_18343_),
    .C(_05476_),
    .Y(_05955_));
 sky130_fd_sc_hd__o22a_2 _34106_ (.A1(_04504_),
    .A2(_18114_),
    .B1(_18343_),
    .B2(_03389_),
    .X(_05956_));
 sky130_fd_sc_hd__nor2_2 _34107_ (.A(_05955_),
    .B(_05956_),
    .Y(_05957_));
 sky130_fd_sc_hd__nand2_2 _34108_ (.A(_00633_),
    .B(_04469_),
    .Y(_05958_));
 sky130_fd_sc_hd__xor2_2 _34109_ (.A(_05957_),
    .B(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__xnor2_2 _34110_ (.A(_05954_),
    .B(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__xnor2_2 _34111_ (.A(_05953_),
    .B(_05960_),
    .Y(_05961_));
 sky130_fd_sc_hd__xnor2_2 _34112_ (.A(_05951_),
    .B(_05961_),
    .Y(_05962_));
 sky130_fd_sc_hd__xnor2_2 _34113_ (.A(_05950_),
    .B(_05962_),
    .Y(_05964_));
 sky130_fd_sc_hd__or2b_2 _34114_ (.A(_05482_),
    .B_N(_05471_),
    .X(_05965_));
 sky130_fd_sc_hd__or2b_2 _34115_ (.A(_05483_),
    .B_N(_05469_),
    .X(_05966_));
 sky130_fd_sc_hd__and2_2 _34116_ (.A(_05965_),
    .B(_05966_),
    .X(_05967_));
 sky130_fd_sc_hd__xor2_2 _34117_ (.A(_05964_),
    .B(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__xnor2_2 _34118_ (.A(_05948_),
    .B(_05968_),
    .Y(_05969_));
 sky130_fd_sc_hd__xor2_2 _34119_ (.A(_05926_),
    .B(_05969_),
    .X(_05970_));
 sky130_fd_sc_hd__xor2_2 _34120_ (.A(_05923_),
    .B(_05970_),
    .X(_05971_));
 sky130_fd_sc_hd__nor2_2 _34121_ (.A(_05527_),
    .B(_05528_),
    .Y(_05972_));
 sky130_fd_sc_hd__a21oi_2 _34122_ (.A1(_05514_),
    .A2(_05529_),
    .B1(_05972_),
    .Y(_05973_));
 sky130_fd_sc_hd__or2b_2 _34123_ (.A(_05556_),
    .B_N(_05559_),
    .X(_05975_));
 sky130_fd_sc_hd__nand2_2 _34124_ (.A(_02984_),
    .B(_18209_),
    .Y(_05976_));
 sky130_fd_sc_hd__nor2_2 _34125_ (.A(_05495_),
    .B(_05976_),
    .Y(_05977_));
 sky130_fd_sc_hd__buf_1 _34126_ (.A(_17409_),
    .X(_05978_));
 sky130_fd_sc_hd__buf_1 _34127_ (.A(_18200_),
    .X(_05979_));
 sky130_fd_sc_hd__buf_1 _34128_ (.A(_18363_),
    .X(_05980_));
 sky130_fd_sc_hd__o22a_2 _34129_ (.A1(_04501_),
    .A2(_05978_),
    .B1(_05979_),
    .B2(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__nor2_2 _34130_ (.A(_05977_),
    .B(_05981_),
    .Y(_05982_));
 sky130_fd_sc_hd__buf_1 _34131_ (.A(_00649_),
    .X(_05983_));
 sky130_fd_sc_hd__nor2_2 _34132_ (.A(_05983_),
    .B(_05500_),
    .Y(_05984_));
 sky130_fd_sc_hd__xnor2_2 _34133_ (.A(_05982_),
    .B(_05984_),
    .Y(_05986_));
 sky130_fd_sc_hd__nor2_2 _34134_ (.A(_16606_),
    .B(_05522_),
    .Y(_05987_));
 sky130_fd_sc_hd__o22a_2 _34135_ (.A1(_16258_),
    .A2(_01066_),
    .B1(_00271_),
    .B2(_00996_),
    .X(_05988_));
 sky130_fd_sc_hd__a21o_2 _34136_ (.A1(_05505_),
    .A2(_05987_),
    .B1(_05988_),
    .X(_05989_));
 sky130_fd_sc_hd__nor2_2 _34137_ (.A(_04847_),
    .B(_04862_),
    .Y(_05990_));
 sky130_fd_sc_hd__xor2_2 _34138_ (.A(_05989_),
    .B(_05990_),
    .X(_05991_));
 sky130_fd_sc_hd__o2bb2ai_2 _34139_ (.A1_N(_05173_),
    .A2_N(_05505_),
    .B1(_05506_),
    .B2(_05508_),
    .Y(_05992_));
 sky130_fd_sc_hd__or2b_2 _34140_ (.A(_05991_),
    .B_N(_05992_),
    .X(_05993_));
 sky130_fd_sc_hd__or2b_2 _34141_ (.A(_05992_),
    .B_N(_05991_),
    .X(_05994_));
 sky130_fd_sc_hd__nand2_2 _34142_ (.A(_05993_),
    .B(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__xor2_2 _34143_ (.A(_05986_),
    .B(_05995_),
    .X(_05997_));
 sky130_fd_sc_hd__a21bo_2 _34144_ (.A1(_05519_),
    .A2(_05523_),
    .B1_N(_05518_),
    .X(_05998_));
 sky130_fd_sc_hd__or3_2 _34145_ (.A(_14949_),
    .B(_01866_),
    .C(_05517_),
    .X(_05999_));
 sky130_fd_sc_hd__o21ai_2 _34146_ (.A1(_14949_),
    .A2(_01866_),
    .B1(_05517_),
    .Y(_06000_));
 sky130_fd_sc_hd__nand2_2 _34147_ (.A(_05999_),
    .B(_06000_),
    .Y(_06001_));
 sky130_fd_sc_hd__nor2_2 _34148_ (.A(_03388_),
    .B(_04162_),
    .Y(_06002_));
 sky130_fd_sc_hd__xnor2_2 _34149_ (.A(_06001_),
    .B(_06002_),
    .Y(_06003_));
 sky130_fd_sc_hd__o21a_2 _34150_ (.A1(_05539_),
    .A2(_05542_),
    .B1(_06003_),
    .X(_06004_));
 sky130_fd_sc_hd__nor3_2 _34151_ (.A(_05539_),
    .B(_05542_),
    .C(_06003_),
    .Y(_06005_));
 sky130_fd_sc_hd__or2_2 _34152_ (.A(_06004_),
    .B(_06005_),
    .X(_06006_));
 sky130_fd_sc_hd__xor2_2 _34153_ (.A(_05998_),
    .B(_06006_),
    .X(_06008_));
 sky130_fd_sc_hd__a21oi_2 _34154_ (.A1(_05222_),
    .A2(_05226_),
    .B1(_05525_),
    .Y(_06009_));
 sky130_fd_sc_hd__a21oi_2 _34155_ (.A1(_05515_),
    .A2(_05526_),
    .B1(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__xor2_2 _34156_ (.A(_06008_),
    .B(_06010_),
    .X(_06011_));
 sky130_fd_sc_hd__xnor2_2 _34157_ (.A(_05997_),
    .B(_06011_),
    .Y(_06012_));
 sky130_fd_sc_hd__xnor2_2 _34158_ (.A(_05975_),
    .B(_06012_),
    .Y(_06013_));
 sky130_fd_sc_hd__or2_2 _34159_ (.A(_05973_),
    .B(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__nand2_2 _34160_ (.A(_05973_),
    .B(_06013_),
    .Y(_06015_));
 sky130_fd_sc_hd__nand2_2 _34161_ (.A(_06014_),
    .B(_06015_),
    .Y(_06016_));
 sky130_fd_sc_hd__or3_2 _34162_ (.A(_02613_),
    .B(_05550_),
    .C(_05233_),
    .X(_06017_));
 sky130_fd_sc_hd__or4_2 _34163_ (.A(_02608_),
    .B(_01605_),
    .C(_02391_),
    .D(_02643_),
    .X(_06019_));
 sky130_fd_sc_hd__a22o_2 _34164_ (.A1(_14593_),
    .A2(_03994_),
    .B1(_03457_),
    .B2(_01039_),
    .X(_06020_));
 sky130_fd_sc_hd__nand2_2 _34165_ (.A(_06019_),
    .B(_06020_),
    .Y(_06021_));
 sky130_fd_sc_hd__or3_2 _34166_ (.A(_01028_),
    .B(_04187_),
    .C(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__buf_1 _34167_ (.A(_04187_),
    .X(_06023_));
 sky130_fd_sc_hd__o21ai_2 _34168_ (.A1(_01028_),
    .A2(_06023_),
    .B1(_06021_),
    .Y(_06024_));
 sky130_fd_sc_hd__and2_2 _34169_ (.A(_06022_),
    .B(_06024_),
    .X(_06025_));
 sky130_fd_sc_hd__xor2_2 _34170_ (.A(_06017_),
    .B(_06025_),
    .X(_06026_));
 sky130_fd_sc_hd__a21oi_2 _34171_ (.A1(_05545_),
    .A2(_05555_),
    .B1(_05553_),
    .Y(_06027_));
 sky130_fd_sc_hd__or2_2 _34172_ (.A(_06026_),
    .B(_06027_),
    .X(_06028_));
 sky130_fd_sc_hd__nand2_2 _34173_ (.A(_06026_),
    .B(_06027_),
    .Y(_06030_));
 sky130_fd_sc_hd__and2_2 _34174_ (.A(_06028_),
    .B(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__a21oi_2 _34175_ (.A1(_05209_),
    .A2(_05215_),
    .B1(_05536_),
    .Y(_06032_));
 sky130_fd_sc_hd__nand2_2 _34176_ (.A(_15641_),
    .B(_05533_),
    .Y(_06033_));
 sky130_fd_sc_hd__o22a_2 _34177_ (.A1(_16288_),
    .A2(_04181_),
    .B1(_04901_),
    .B2(_18791_),
    .X(_06034_));
 sky130_fd_sc_hd__a31o_2 _34178_ (.A1(_01785_),
    .A2(_13544_),
    .A3(_03064_),
    .B1(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__nand2_2 _34179_ (.A(_06033_),
    .B(_06035_),
    .Y(_06036_));
 sky130_fd_sc_hd__or2_2 _34180_ (.A(_06033_),
    .B(_06035_),
    .X(_06037_));
 sky130_fd_sc_hd__or2_2 _34181_ (.A(_05536_),
    .B(_06035_),
    .X(_06038_));
 sky130_fd_sc_hd__a21o_2 _34182_ (.A1(_05209_),
    .A2(_05215_),
    .B1(_06038_),
    .X(_06039_));
 sky130_fd_sc_hd__o211a_2 _34183_ (.A1(_06032_),
    .A2(_06036_),
    .B1(_06037_),
    .C1(_06039_),
    .X(_06041_));
 sky130_fd_sc_hd__xnor2_2 _34184_ (.A(_06031_),
    .B(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__xor2_2 _34185_ (.A(_05561_),
    .B(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__xnor2_2 _34186_ (.A(_06016_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__a21oi_2 _34187_ (.A1(_05532_),
    .A2(_05566_),
    .B1(_05564_),
    .Y(_06045_));
 sky130_fd_sc_hd__xnor2_2 _34188_ (.A(_06044_),
    .B(_06045_),
    .Y(_06046_));
 sky130_fd_sc_hd__xnor2_2 _34189_ (.A(_05971_),
    .B(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__or2_2 _34190_ (.A(_05567_),
    .B(_05570_),
    .X(_06048_));
 sky130_fd_sc_hd__o21a_2 _34191_ (.A1(_05490_),
    .A2(_05571_),
    .B1(_06048_),
    .X(_06049_));
 sky130_fd_sc_hd__xnor2_2 _34192_ (.A(_06047_),
    .B(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__xnor2_2 _34193_ (.A(_05922_),
    .B(_06050_),
    .Y(_06052_));
 sky130_fd_sc_hd__or2b_2 _34194_ (.A(_05574_),
    .B_N(_05572_),
    .X(_06053_));
 sky130_fd_sc_hd__a21boi_2 _34195_ (.A1(_05433_),
    .A2(_05575_),
    .B1_N(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__nor2_2 _34196_ (.A(_06052_),
    .B(_06054_),
    .Y(_06055_));
 sky130_fd_sc_hd__nand2_2 _34197_ (.A(_06052_),
    .B(_06054_),
    .Y(_06056_));
 sky130_fd_sc_hd__and2b_2 _34198_ (.A_N(_06055_),
    .B(_06056_),
    .X(_06057_));
 sky130_fd_sc_hd__xnor2_2 _34199_ (.A(_05913_),
    .B(_06057_),
    .Y(_06058_));
 sky130_fd_sc_hd__a21o_2 _34200_ (.A1(_05116_),
    .A2(_05582_),
    .B1(_05580_),
    .X(_06059_));
 sky130_fd_sc_hd__xnor2_2 _34201_ (.A(_06058_),
    .B(_06059_),
    .Y(_06060_));
 sky130_fd_sc_hd__nor2_2 _34202_ (.A(_05586_),
    .B(_05589_),
    .Y(_06061_));
 sky130_fd_sc_hd__xnor2_2 _34203_ (.A(_06060_),
    .B(_06061_),
    .Y(_06063_));
 sky130_fd_sc_hd__xnor2_2 _34204_ (.A(_05912_),
    .B(_06063_),
    .Y(_06064_));
 sky130_fd_sc_hd__xnor2_2 _34205_ (.A(_13489_),
    .B(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__o31a_2 _34206_ (.A1(_05589_),
    .A2(_05591_),
    .A3(_05751_),
    .B1(_05753_),
    .X(_06066_));
 sky130_fd_sc_hd__xor2_2 _34207_ (.A(_06065_),
    .B(_06066_),
    .X(_06067_));
 sky130_fd_sc_hd__nor2_2 _34208_ (.A(_05756_),
    .B(_05757_),
    .Y(_06068_));
 sky130_fd_sc_hd__and2b_2 _34209_ (.A_N(_05767_),
    .B(_05758_),
    .X(_06069_));
 sky130_fd_sc_hd__nor2_2 _34210_ (.A(_06068_),
    .B(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__xnor2_2 _34211_ (.A(_06067_),
    .B(_06070_),
    .Y(_06071_));
 sky130_fd_sc_hd__and2_2 _34212_ (.A(_13616_),
    .B(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__or2_2 _34213_ (.A(_13616_),
    .B(_06071_),
    .X(_06074_));
 sky130_fd_sc_hd__and2b_2 _34214_ (.A_N(_06072_),
    .B(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__and2b_2 _34215_ (.A_N(_05782_),
    .B(_05771_),
    .X(_06076_));
 sky130_fd_sc_hd__nor2_2 _34216_ (.A(_05769_),
    .B(_06076_),
    .Y(_06077_));
 sky130_fd_sc_hd__xnor2_2 _34217_ (.A(_06075_),
    .B(_06077_),
    .Y(oO[73]));
 sky130_fd_sc_hd__a21o_2 _34218_ (.A1(_05769_),
    .A2(_06074_),
    .B1(_06072_),
    .X(_06078_));
 sky130_fd_sc_hd__a21oi_2 _34219_ (.A1(_06076_),
    .A2(_06075_),
    .B1(_06078_),
    .Y(_06079_));
 sky130_fd_sc_hd__or2b_2 _34220_ (.A(_05912_),
    .B_N(_06063_),
    .X(_06080_));
 sky130_fd_sc_hd__nand2_2 _34221_ (.A(_13489_),
    .B(_06064_),
    .Y(_06081_));
 sky130_fd_sc_hd__inv_2 _34222_ (.A(_13768_),
    .Y(_06082_));
 sky130_fd_sc_hd__or2b_2 _34223_ (.A(_05969_),
    .B_N(_05926_),
    .X(_06084_));
 sky130_fd_sc_hd__or2b_2 _34224_ (.A(_05970_),
    .B_N(_05923_),
    .X(_06085_));
 sky130_fd_sc_hd__and2b_2 _34225_ (.A_N(_05945_),
    .B(_05946_),
    .X(_06086_));
 sky130_fd_sc_hd__and2b_2 _34226_ (.A_N(_05927_),
    .B(_05947_),
    .X(_06087_));
 sky130_fd_sc_hd__nor2_2 _34227_ (.A(_06086_),
    .B(_06087_),
    .Y(_06088_));
 sky130_fd_sc_hd__a21oi_2 _34228_ (.A1(_06084_),
    .A2(_06085_),
    .B1(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__and3_2 _34229_ (.A(_06084_),
    .B(_06085_),
    .C(_06088_),
    .X(_06090_));
 sky130_fd_sc_hd__nor2_2 _34230_ (.A(_06089_),
    .B(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__nor2_2 _34231_ (.A(_05964_),
    .B(_05967_),
    .Y(_06092_));
 sky130_fd_sc_hd__a21o_2 _34232_ (.A1(_05948_),
    .A2(_05968_),
    .B1(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__o21ai_2 _34233_ (.A1(_05975_),
    .A2(_06012_),
    .B1(_06014_),
    .Y(_06095_));
 sky130_fd_sc_hd__o31ai_2 _34234_ (.A1(_01797_),
    .A2(_05441_),
    .A3(_05933_),
    .B1(_05929_),
    .Y(_06096_));
 sky130_fd_sc_hd__or3_2 _34235_ (.A(_02463_),
    .B(_02317_),
    .C(_05928_),
    .X(_06097_));
 sky130_fd_sc_hd__a2bb2o_2 _34236_ (.A1_N(_01583_),
    .A2_N(_02317_),
    .B1(_02928_),
    .B2(_02983_),
    .X(_06098_));
 sky130_fd_sc_hd__nand2_2 _34237_ (.A(_06097_),
    .B(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__nor2_2 _34238_ (.A(_01576_),
    .B(_03318_),
    .Y(_06100_));
 sky130_fd_sc_hd__xnor2_2 _34239_ (.A(_06099_),
    .B(_06100_),
    .Y(_06101_));
 sky130_fd_sc_hd__nand2_2 _34240_ (.A(_00633_),
    .B(_00566_),
    .Y(_06102_));
 sky130_fd_sc_hd__o22a_2 _34241_ (.A1(_01832_),
    .A2(_02940_),
    .B1(_02311_),
    .B2(_03378_),
    .X(_06103_));
 sky130_fd_sc_hd__o21bai_2 _34242_ (.A1(_05936_),
    .A2(_06102_),
    .B1_N(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__nand2_2 _34243_ (.A(_02994_),
    .B(_03327_),
    .Y(_06106_));
 sky130_fd_sc_hd__xnor2_2 _34244_ (.A(_06104_),
    .B(_06106_),
    .Y(_06107_));
 sky130_fd_sc_hd__or2_2 _34245_ (.A(_05452_),
    .B(_05936_),
    .X(_06108_));
 sky130_fd_sc_hd__o21a_2 _34246_ (.A1(_05937_),
    .A2(_05938_),
    .B1(_06108_),
    .X(_06109_));
 sky130_fd_sc_hd__or2_2 _34247_ (.A(_06107_),
    .B(_06109_),
    .X(_06110_));
 sky130_fd_sc_hd__nand2_2 _34248_ (.A(_06107_),
    .B(_06109_),
    .Y(_06111_));
 sky130_fd_sc_hd__and2_2 _34249_ (.A(_06110_),
    .B(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__nand2_2 _34250_ (.A(_06101_),
    .B(_06112_),
    .Y(_06113_));
 sky130_fd_sc_hd__or2_2 _34251_ (.A(_06101_),
    .B(_06112_),
    .X(_06114_));
 sky130_fd_sc_hd__nand2_2 _34252_ (.A(_06113_),
    .B(_06114_),
    .Y(_06115_));
 sky130_fd_sc_hd__a21o_2 _34253_ (.A1(_05935_),
    .A2(_05944_),
    .B1(_05942_),
    .X(_06117_));
 sky130_fd_sc_hd__xnor2_2 _34254_ (.A(_06115_),
    .B(_06117_),
    .Y(_06118_));
 sky130_fd_sc_hd__xnor2_2 _34255_ (.A(_06096_),
    .B(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__or2b_2 _34256_ (.A(_05959_),
    .B_N(_05954_),
    .X(_06120_));
 sky130_fd_sc_hd__a21bo_2 _34257_ (.A1(_05953_),
    .A2(_05960_),
    .B1_N(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__o21a_2 _34258_ (.A1(_05986_),
    .A2(_05995_),
    .B1(_05993_),
    .X(_06122_));
 sky130_fd_sc_hd__a31o_2 _34259_ (.A1(_00633_),
    .A2(_04469_),
    .A3(_05957_),
    .B1(_05955_),
    .X(_06123_));
 sky130_fd_sc_hd__a31o_2 _34260_ (.A1(_01837_),
    .A2(_03345_),
    .A3(_05982_),
    .B1(_05977_),
    .X(_06124_));
 sky130_fd_sc_hd__and4_2 _34261_ (.A(_04837_),
    .B(_01837_),
    .C(_18328_),
    .D(_18734_),
    .X(_06125_));
 sky130_fd_sc_hd__o22a_2 _34262_ (.A1(_00649_),
    .A2(_18114_),
    .B1(_18343_),
    .B2(_04504_),
    .X(_06126_));
 sky130_fd_sc_hd__nor2_2 _34263_ (.A(_06125_),
    .B(_06126_),
    .Y(_06128_));
 sky130_fd_sc_hd__nand2_2 _34264_ (.A(_01040_),
    .B(_02956_),
    .Y(_06129_));
 sky130_fd_sc_hd__xor2_2 _34265_ (.A(_06128_),
    .B(_06129_),
    .X(_06130_));
 sky130_fd_sc_hd__xnor2_2 _34266_ (.A(_06124_),
    .B(_06130_),
    .Y(_06131_));
 sky130_fd_sc_hd__xnor2_2 _34267_ (.A(_06123_),
    .B(_06131_),
    .Y(_06132_));
 sky130_fd_sc_hd__xnor2_2 _34268_ (.A(_06122_),
    .B(_06132_),
    .Y(_06133_));
 sky130_fd_sc_hd__xnor2_2 _34269_ (.A(_06121_),
    .B(_06133_),
    .Y(_06134_));
 sky130_fd_sc_hd__nor2_2 _34270_ (.A(_05951_),
    .B(_05961_),
    .Y(_06135_));
 sky130_fd_sc_hd__nor2_2 _34271_ (.A(_05950_),
    .B(_05962_),
    .Y(_06136_));
 sky130_fd_sc_hd__nor2_2 _34272_ (.A(_06135_),
    .B(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__xnor2_2 _34273_ (.A(_06134_),
    .B(_06137_),
    .Y(_06139_));
 sky130_fd_sc_hd__xnor2_2 _34274_ (.A(_06119_),
    .B(_06139_),
    .Y(_06140_));
 sky130_fd_sc_hd__xnor2_2 _34275_ (.A(_06095_),
    .B(_06140_),
    .Y(_06141_));
 sky130_fd_sc_hd__xor2_2 _34276_ (.A(_06093_),
    .B(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__and2_2 _34277_ (.A(_06031_),
    .B(_06041_),
    .X(_06143_));
 sky130_fd_sc_hd__o22a_2 _34278_ (.A1(_01797_),
    .A2(_04181_),
    .B1(_04901_),
    .B2(_02613_),
    .X(_06144_));
 sky130_fd_sc_hd__a31o_2 _34279_ (.A1(_00999_),
    .A2(_13889_),
    .A3(_05533_),
    .B1(_06144_),
    .X(_06145_));
 sky130_fd_sc_hd__o21a_2 _34280_ (.A1(_16275_),
    .A2(_03068_),
    .B1(_06037_),
    .X(_06146_));
 sky130_fd_sc_hd__and2_2 _34281_ (.A(_06039_),
    .B(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__xor2_2 _34282_ (.A(_06145_),
    .B(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__nand2_2 _34283_ (.A(_14593_),
    .B(_03457_),
    .Y(_06150_));
 sky130_fd_sc_hd__nor2_2 _34284_ (.A(_02608_),
    .B(_02652_),
    .Y(_06151_));
 sky130_fd_sc_hd__xnor2_2 _34285_ (.A(_06150_),
    .B(_06151_),
    .Y(_06152_));
 sky130_fd_sc_hd__and3_2 _34286_ (.A(_03023_),
    .B(_03994_),
    .C(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__buf_1 _34287_ (.A(_03994_),
    .X(_06154_));
 sky130_fd_sc_hd__a21oi_2 _34288_ (.A1(_03023_),
    .A2(_06154_),
    .B1(_06152_),
    .Y(_06155_));
 sky130_fd_sc_hd__o211ai_2 _34289_ (.A1(_05233_),
    .A2(_06025_),
    .B1(_13889_),
    .C1(_04905_),
    .Y(_06156_));
 sky130_fd_sc_hd__or3_2 _34290_ (.A(_06153_),
    .B(_06155_),
    .C(_06156_),
    .X(_06157_));
 sky130_fd_sc_hd__o21ai_2 _34291_ (.A1(_06153_),
    .A2(_06155_),
    .B1(_06156_),
    .Y(_06158_));
 sky130_fd_sc_hd__and2_2 _34292_ (.A(_06157_),
    .B(_06158_),
    .X(_06159_));
 sky130_fd_sc_hd__xor2_2 _34293_ (.A(_06148_),
    .B(_06159_),
    .X(_06161_));
 sky130_fd_sc_hd__xnor2_2 _34294_ (.A(_06143_),
    .B(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__nor2_2 _34295_ (.A(_06008_),
    .B(_06010_),
    .Y(_06163_));
 sky130_fd_sc_hd__a21o_2 _34296_ (.A1(_05997_),
    .A2(_06011_),
    .B1(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__or2_2 _34297_ (.A(_05980_),
    .B(_04862_),
    .X(_06165_));
 sky130_fd_sc_hd__xor2_2 _34298_ (.A(_05976_),
    .B(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__nor2_2 _34299_ (.A(_04501_),
    .B(_05500_),
    .Y(_06167_));
 sky130_fd_sc_hd__xnor2_2 _34300_ (.A(_06166_),
    .B(_06167_),
    .Y(_06168_));
 sky130_fd_sc_hd__nor2_2 _34301_ (.A(_00996_),
    .B(_04162_),
    .Y(_06169_));
 sky130_fd_sc_hd__nand2_2 _34302_ (.A(_05987_),
    .B(_06169_),
    .Y(_06170_));
 sky130_fd_sc_hd__or2_2 _34303_ (.A(_05987_),
    .B(_06169_),
    .X(_06172_));
 sky130_fd_sc_hd__and2_2 _34304_ (.A(_06170_),
    .B(_06172_),
    .X(_06173_));
 sky130_fd_sc_hd__nor2_2 _34305_ (.A(_04847_),
    .B(_05504_),
    .Y(_06174_));
 sky130_fd_sc_hd__xnor2_2 _34306_ (.A(_06173_),
    .B(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__inv_2 _34307_ (.A(_05989_),
    .Y(_06176_));
 sky130_fd_sc_hd__a22o_2 _34308_ (.A1(_05505_),
    .A2(_05987_),
    .B1(_06176_),
    .B2(_05990_),
    .X(_06177_));
 sky130_fd_sc_hd__or2b_2 _34309_ (.A(_06175_),
    .B_N(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__or2b_2 _34310_ (.A(_06177_),
    .B_N(_06175_),
    .X(_06179_));
 sky130_fd_sc_hd__nand2_2 _34311_ (.A(_06178_),
    .B(_06179_),
    .Y(_06180_));
 sky130_fd_sc_hd__xor2_2 _34312_ (.A(_06168_),
    .B(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__and2b_2 _34313_ (.A_N(_06006_),
    .B(_05998_),
    .X(_06183_));
 sky130_fd_sc_hd__a21bo_2 _34314_ (.A1(_06000_),
    .A2(_06002_),
    .B1_N(_05999_),
    .X(_06184_));
 sky130_fd_sc_hd__nor2_2 _34315_ (.A(_15155_),
    .B(_02647_),
    .Y(_06185_));
 sky130_fd_sc_hd__and3_2 _34316_ (.A(_01033_),
    .B(_03438_),
    .C(_06185_),
    .X(_06186_));
 sky130_fd_sc_hd__o22a_2 _34317_ (.A1(_15155_),
    .A2(_01866_),
    .B1(_04187_),
    .B2(_14949_),
    .X(_06187_));
 sky130_fd_sc_hd__nor2_2 _34318_ (.A(_06186_),
    .B(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__nor2_2 _34319_ (.A(_03388_),
    .B(_01070_),
    .Y(_06189_));
 sky130_fd_sc_hd__xnor2_2 _34320_ (.A(_06188_),
    .B(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__a21o_2 _34321_ (.A1(_06019_),
    .A2(_06022_),
    .B1(_06190_),
    .X(_06191_));
 sky130_fd_sc_hd__nand3_2 _34322_ (.A(_06019_),
    .B(_06022_),
    .C(_06190_),
    .Y(_06192_));
 sky130_fd_sc_hd__nand2_2 _34323_ (.A(_06191_),
    .B(_06192_),
    .Y(_06194_));
 sky130_fd_sc_hd__xnor2_2 _34324_ (.A(_06184_),
    .B(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__o21a_2 _34325_ (.A1(_06004_),
    .A2(_06183_),
    .B1(_06195_),
    .X(_06196_));
 sky130_fd_sc_hd__nor3_2 _34326_ (.A(_06004_),
    .B(_06183_),
    .C(_06195_),
    .Y(_06197_));
 sky130_fd_sc_hd__nor2_2 _34327_ (.A(_06196_),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__xnor2_2 _34328_ (.A(_06181_),
    .B(_06198_),
    .Y(_06199_));
 sky130_fd_sc_hd__nor2_2 _34329_ (.A(_06028_),
    .B(_06199_),
    .Y(_06200_));
 sky130_fd_sc_hd__and2_2 _34330_ (.A(_06028_),
    .B(_06199_),
    .X(_06201_));
 sky130_fd_sc_hd__nor2_2 _34331_ (.A(_06200_),
    .B(_06201_),
    .Y(_06202_));
 sky130_fd_sc_hd__xnor2_2 _34332_ (.A(_06164_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__xor2_2 _34333_ (.A(_06162_),
    .B(_06203_),
    .X(_06205_));
 sky130_fd_sc_hd__nor2_2 _34334_ (.A(_05561_),
    .B(_06042_),
    .Y(_06206_));
 sky130_fd_sc_hd__a31o_2 _34335_ (.A1(_06014_),
    .A2(_06015_),
    .A3(_06043_),
    .B1(_06206_),
    .X(_06207_));
 sky130_fd_sc_hd__xnor2_2 _34336_ (.A(_06205_),
    .B(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__xnor2_2 _34337_ (.A(_06142_),
    .B(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__and2b_2 _34338_ (.A_N(_06044_),
    .B(_06045_),
    .X(_06210_));
 sky130_fd_sc_hd__or2b_2 _34339_ (.A(_06045_),
    .B_N(_06044_),
    .X(_06211_));
 sky130_fd_sc_hd__o21ai_2 _34340_ (.A1(_05971_),
    .A2(_06210_),
    .B1(_06211_),
    .Y(_06212_));
 sky130_fd_sc_hd__xnor2_2 _34341_ (.A(_06209_),
    .B(_06212_),
    .Y(_06213_));
 sky130_fd_sc_hd__xnor2_2 _34342_ (.A(_06091_),
    .B(_06213_),
    .Y(_06214_));
 sky130_fd_sc_hd__and2b_2 _34343_ (.A_N(_06049_),
    .B(_06047_),
    .X(_06216_));
 sky130_fd_sc_hd__a21o_2 _34344_ (.A1(_05922_),
    .A2(_06050_),
    .B1(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__xnor2_2 _34345_ (.A(_06214_),
    .B(_06217_),
    .Y(_06218_));
 sky130_fd_sc_hd__xnor2_2 _34346_ (.A(_05920_),
    .B(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__a21oi_2 _34347_ (.A1(_05913_),
    .A2(_06056_),
    .B1(_06055_),
    .Y(_06220_));
 sky130_fd_sc_hd__xnor2_2 _34348_ (.A(_06219_),
    .B(_06220_),
    .Y(_06221_));
 sky130_fd_sc_hd__or2b_2 _34349_ (.A(_06059_),
    .B_N(_06058_),
    .X(_06222_));
 sky130_fd_sc_hd__and2b_2 _34350_ (.A_N(_06058_),
    .B(_06059_),
    .X(_06223_));
 sky130_fd_sc_hd__a21oi_2 _34351_ (.A1(_05586_),
    .A2(_06222_),
    .B1(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__a21boi_2 _34352_ (.A1(_05589_),
    .A2(_06060_),
    .B1_N(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__xnor2_2 _34353_ (.A(_06221_),
    .B(_06225_),
    .Y(_06227_));
 sky130_fd_sc_hd__and3b_2 _34354_ (.A_N(_05274_),
    .B(iX[63]),
    .C(iY[43]),
    .X(_06228_));
 sky130_fd_sc_hd__and2_2 _34355_ (.A(iY[45]),
    .B(iX[62]),
    .X(_06229_));
 sky130_fd_sc_hd__and3_2 _34356_ (.A(iY[44]),
    .B(iX[61]),
    .C(_06229_),
    .X(_06230_));
 sky130_fd_sc_hd__a22oi_2 _34357_ (.A1(iY[45]),
    .A2(iX[61]),
    .B1(iX[62]),
    .B2(iY[44]),
    .Y(_06231_));
 sky130_fd_sc_hd__nor2_2 _34358_ (.A(_06230_),
    .B(_06231_),
    .Y(_06232_));
 sky130_fd_sc_hd__a21oi_2 _34359_ (.A1(iY[46]),
    .A2(iX[60]),
    .B1(_06232_),
    .Y(_06233_));
 sky130_fd_sc_hd__and3_2 _34360_ (.A(iY[46]),
    .B(iX[60]),
    .C(_06232_),
    .X(_06234_));
 sky130_fd_sc_hd__nor2_2 _34361_ (.A(_06233_),
    .B(_06234_),
    .Y(_06235_));
 sky130_fd_sc_hd__xnor2_2 _34362_ (.A(_06228_),
    .B(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__or2b_2 _34363_ (.A(_05786_),
    .B_N(_05788_),
    .X(_06238_));
 sky130_fd_sc_hd__a21bo_2 _34364_ (.A1(_05789_),
    .A2(_05794_),
    .B1_N(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__xor2_2 _34365_ (.A(_06236_),
    .B(_06239_),
    .X(_06240_));
 sky130_fd_sc_hd__a21o_2 _34366_ (.A1(_05818_),
    .A2(_05660_),
    .B1(_05830_),
    .X(_06241_));
 sky130_fd_sc_hd__and4_2 _34367_ (.A(iX[52]),
    .B(iX[53]),
    .C(iY[53]),
    .D(iY[54]),
    .X(_06242_));
 sky130_fd_sc_hd__a22oi_2 _34368_ (.A1(iX[53]),
    .A2(iY[53]),
    .B1(iY[54]),
    .B2(iX[52]),
    .Y(_06243_));
 sky130_fd_sc_hd__nor2_2 _34369_ (.A(_06242_),
    .B(_06243_),
    .Y(_06244_));
 sky130_fd_sc_hd__nand2_2 _34370_ (.A(iX[51]),
    .B(iY[55]),
    .Y(_06245_));
 sky130_fd_sc_hd__xnor2_2 _34371_ (.A(_06244_),
    .B(_06245_),
    .Y(_06246_));
 sky130_fd_sc_hd__and4_2 _34372_ (.A(iY[50]),
    .B(iY[51]),
    .C(iX[55]),
    .D(iX[56]),
    .X(_06247_));
 sky130_fd_sc_hd__a22oi_2 _34373_ (.A1(iY[51]),
    .A2(iX[55]),
    .B1(iX[56]),
    .B2(iY[50]),
    .Y(_06249_));
 sky130_fd_sc_hd__nor2_2 _34374_ (.A(_06247_),
    .B(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__nand2_2 _34375_ (.A(iY[52]),
    .B(iX[54]),
    .Y(_06251_));
 sky130_fd_sc_hd__xnor2_2 _34376_ (.A(_06250_),
    .B(_06251_),
    .Y(_06252_));
 sky130_fd_sc_hd__o21ba_2 _34377_ (.A1(_05808_),
    .A2(_05811_),
    .B1_N(_05807_),
    .X(_06253_));
 sky130_fd_sc_hd__xnor2_2 _34378_ (.A(_06252_),
    .B(_06253_),
    .Y(_06254_));
 sky130_fd_sc_hd__and2_2 _34379_ (.A(_06246_),
    .B(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__nor2_2 _34380_ (.A(_06246_),
    .B(_06254_),
    .Y(_06256_));
 sky130_fd_sc_hd__or2_2 _34381_ (.A(_06255_),
    .B(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__nand2_2 _34382_ (.A(_05819_),
    .B(_05829_),
    .Y(_06258_));
 sky130_fd_sc_hd__o21ba_2 _34383_ (.A1(_05791_),
    .A2(_05793_),
    .B1_N(_05790_),
    .X(_06260_));
 sky130_fd_sc_hd__and4_2 _34384_ (.A(iY[47]),
    .B(iY[48]),
    .C(iX[58]),
    .D(iX[59]),
    .X(_06261_));
 sky130_fd_sc_hd__a22oi_2 _34385_ (.A1(iY[48]),
    .A2(iX[58]),
    .B1(iX[59]),
    .B2(iY[47]),
    .Y(_06262_));
 sky130_fd_sc_hd__nor2_2 _34386_ (.A(_06261_),
    .B(_06262_),
    .Y(_06263_));
 sky130_fd_sc_hd__nand2_2 _34387_ (.A(iY[49]),
    .B(iX[57]),
    .Y(_06264_));
 sky130_fd_sc_hd__xnor2_2 _34388_ (.A(_06263_),
    .B(_06264_),
    .Y(_06265_));
 sky130_fd_sc_hd__xnor2_2 _34389_ (.A(_06260_),
    .B(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__o21ai_2 _34390_ (.A1(_05821_),
    .A2(_05825_),
    .B1(_06266_),
    .Y(_06267_));
 sky130_fd_sc_hd__or3_2 _34391_ (.A(_05821_),
    .B(_05825_),
    .C(_06266_),
    .X(_06268_));
 sky130_fd_sc_hd__nand2_2 _34392_ (.A(_06267_),
    .B(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__a21oi_2 _34393_ (.A1(_05827_),
    .A2(_06258_),
    .B1(_06269_),
    .Y(_06271_));
 sky130_fd_sc_hd__and3_2 _34394_ (.A(_05827_),
    .B(_06258_),
    .C(_06269_),
    .X(_06272_));
 sky130_fd_sc_hd__or3_2 _34395_ (.A(_06257_),
    .B(_06271_),
    .C(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__o21ai_2 _34396_ (.A1(_06271_),
    .A2(_06272_),
    .B1(_06257_),
    .Y(_06274_));
 sky130_fd_sc_hd__and3_2 _34397_ (.A(_05796_),
    .B(_06273_),
    .C(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__a21oi_2 _34398_ (.A1(_06273_),
    .A2(_06274_),
    .B1(_05796_),
    .Y(_06276_));
 sky130_fd_sc_hd__a211oi_2 _34399_ (.A1(_06241_),
    .A2(_05834_),
    .B1(_06275_),
    .C1(_06276_),
    .Y(_06277_));
 sky130_fd_sc_hd__o211a_2 _34400_ (.A1(_06275_),
    .A2(_06276_),
    .B1(_06241_),
    .C1(_05834_),
    .X(_06278_));
 sky130_fd_sc_hd__or3_2 _34401_ (.A(_06240_),
    .B(_06277_),
    .C(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__inv_2 _34402_ (.A(_06279_),
    .Y(_06280_));
 sky130_fd_sc_hd__o21a_2 _34403_ (.A1(_06277_),
    .A2(_06278_),
    .B1(_06240_),
    .X(_06282_));
 sky130_fd_sc_hd__o21ai_2 _34404_ (.A1(_06280_),
    .A2(_06282_),
    .B1(_05840_),
    .Y(_06283_));
 sky130_fd_sc_hd__or3_2 _34405_ (.A(_05840_),
    .B(_06280_),
    .C(_06282_),
    .X(_06284_));
 sky130_fd_sc_hd__inv_2 _34406_ (.A(_05884_),
    .Y(_06285_));
 sky130_fd_sc_hd__and4_2 _34407_ (.A(iX[46]),
    .B(iX[47]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_06286_));
 sky130_fd_sc_hd__a22oi_2 _34408_ (.A1(iX[47]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[46]),
    .Y(_06287_));
 sky130_fd_sc_hd__nor2_2 _34409_ (.A(_06286_),
    .B(_06287_),
    .Y(_06288_));
 sky130_fd_sc_hd__nand2_2 _34410_ (.A(iX[45]),
    .B(iY[61]),
    .Y(_06289_));
 sky130_fd_sc_hd__xnor2_2 _34411_ (.A(_06288_),
    .B(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__o21ba_2 _34412_ (.A1(_05850_),
    .A2(_05852_),
    .B1_N(_05849_),
    .X(_06291_));
 sky130_fd_sc_hd__xnor2_2 _34413_ (.A(_06290_),
    .B(_06291_),
    .Y(_06293_));
 sky130_fd_sc_hd__and2_2 _34414_ (.A(iX[44]),
    .B(iY[62]),
    .X(_06294_));
 sky130_fd_sc_hd__or2_2 _34415_ (.A(_06293_),
    .B(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__nand2_2 _34416_ (.A(_06293_),
    .B(_06294_),
    .Y(_06296_));
 sky130_fd_sc_hd__and2b_2 _34417_ (.A_N(_05855_),
    .B(_05854_),
    .X(_06297_));
 sky130_fd_sc_hd__a31o_2 _34418_ (.A1(iX[43]),
    .A2(iY[62]),
    .A3(_05856_),
    .B1(_06297_),
    .X(_06298_));
 sky130_fd_sc_hd__nand3_2 _34419_ (.A(_06295_),
    .B(_06296_),
    .C(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__a21o_2 _34420_ (.A1(_06295_),
    .A2(_06296_),
    .B1(_06298_),
    .X(_06300_));
 sky130_fd_sc_hd__nand2_2 _34421_ (.A(_06299_),
    .B(_06300_),
    .Y(_06301_));
 sky130_fd_sc_hd__nand2_2 _34422_ (.A(iX[43]),
    .B(iY[63]),
    .Y(_06302_));
 sky130_fd_sc_hd__nand2_2 _34423_ (.A(_06301_),
    .B(_06302_),
    .Y(_06304_));
 sky130_fd_sc_hd__or2_2 _34424_ (.A(_06301_),
    .B(_06302_),
    .X(_06305_));
 sky130_fd_sc_hd__and2_2 _34425_ (.A(_06304_),
    .B(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__or2b_2 _34426_ (.A(_05870_),
    .B_N(_05876_),
    .X(_06307_));
 sky130_fd_sc_hd__or2b_2 _34427_ (.A(_05869_),
    .B_N(_05877_),
    .X(_06308_));
 sky130_fd_sc_hd__and2b_2 _34428_ (.A_N(_05813_),
    .B(_05812_),
    .X(_06309_));
 sky130_fd_sc_hd__o21ba_2 _34429_ (.A1(_05872_),
    .A2(_05874_),
    .B1_N(_05871_),
    .X(_06310_));
 sky130_fd_sc_hd__o21ba_2 _34430_ (.A1(_05803_),
    .A2(_05805_),
    .B1_N(_05802_),
    .X(_06311_));
 sky130_fd_sc_hd__and4_2 _34431_ (.A(iX[49]),
    .B(iX[50]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_06312_));
 sky130_fd_sc_hd__a22oi_2 _34432_ (.A1(iX[50]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[49]),
    .Y(_06313_));
 sky130_fd_sc_hd__nor2_2 _34433_ (.A(_06312_),
    .B(_06313_),
    .Y(_06315_));
 sky130_fd_sc_hd__nand2_2 _34434_ (.A(iX[48]),
    .B(iY[58]),
    .Y(_06316_));
 sky130_fd_sc_hd__xnor2_2 _34435_ (.A(_06315_),
    .B(_06316_),
    .Y(_06317_));
 sky130_fd_sc_hd__xnor2_2 _34436_ (.A(_06311_),
    .B(_06317_),
    .Y(_06318_));
 sky130_fd_sc_hd__xnor2_2 _34437_ (.A(_06310_),
    .B(_06318_),
    .Y(_06319_));
 sky130_fd_sc_hd__o21a_2 _34438_ (.A1(_06309_),
    .A2(_05815_),
    .B1(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__nor3_2 _34439_ (.A(_06309_),
    .B(_05815_),
    .C(_06319_),
    .Y(_06321_));
 sky130_fd_sc_hd__a211oi_2 _34440_ (.A1(_06307_),
    .A2(_06308_),
    .B1(_06320_),
    .C1(_06321_),
    .Y(_06322_));
 sky130_fd_sc_hd__o211a_2 _34441_ (.A1(_06320_),
    .A2(_06321_),
    .B1(_06307_),
    .C1(_06308_),
    .X(_06323_));
 sky130_fd_sc_hd__nor2_2 _34442_ (.A(_05879_),
    .B(_05881_),
    .Y(_06324_));
 sky130_fd_sc_hd__or3_2 _34443_ (.A(_06322_),
    .B(_06323_),
    .C(_06324_),
    .X(_06326_));
 sky130_fd_sc_hd__o21ai_2 _34444_ (.A1(_06322_),
    .A2(_06323_),
    .B1(_06324_),
    .Y(_06327_));
 sky130_fd_sc_hd__and3_2 _34445_ (.A(_06306_),
    .B(_06326_),
    .C(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__a21oi_2 _34446_ (.A1(_06326_),
    .A2(_06327_),
    .B1(_06306_),
    .Y(_06329_));
 sky130_fd_sc_hd__nor2_2 _34447_ (.A(_06328_),
    .B(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__o21ai_2 _34448_ (.A1(_05836_),
    .A2(_05838_),
    .B1(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__or3_2 _34449_ (.A(_05836_),
    .B(_05838_),
    .C(_06330_),
    .X(_06332_));
 sky130_fd_sc_hd__o211ai_2 _34450_ (.A1(_06285_),
    .A2(_05887_),
    .B1(_06331_),
    .C1(_06332_),
    .Y(_06333_));
 sky130_fd_sc_hd__a211o_2 _34451_ (.A1(_06331_),
    .A2(_06332_),
    .B1(_06285_),
    .C1(_05887_),
    .X(_06334_));
 sky130_fd_sc_hd__nand4_2 _34452_ (.A(_06283_),
    .B(_06284_),
    .C(_06333_),
    .D(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__a22o_2 _34453_ (.A1(_06283_),
    .A2(_06284_),
    .B1(_06333_),
    .B2(_06334_),
    .X(_06337_));
 sky130_fd_sc_hd__nand2_2 _34454_ (.A(_05843_),
    .B(_05894_),
    .Y(_06338_));
 sky130_fd_sc_hd__and3_2 _34455_ (.A(_06335_),
    .B(_06337_),
    .C(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__a21oi_2 _34456_ (.A1(_06335_),
    .A2(_06337_),
    .B1(_06338_),
    .Y(_06340_));
 sky130_fd_sc_hd__a211oi_2 _34457_ (.A1(_05889_),
    .A2(_05892_),
    .B1(_06339_),
    .C1(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__o211a_2 _34458_ (.A1(_06339_),
    .A2(_06340_),
    .B1(_05889_),
    .C1(_05892_),
    .X(_06342_));
 sky130_fd_sc_hd__nor2_2 _34459_ (.A(_06341_),
    .B(_06342_),
    .Y(_06343_));
 sky130_fd_sc_hd__o21a_2 _34460_ (.A1(_05898_),
    .A2(_05900_),
    .B1(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__inv_2 _34461_ (.A(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__or3_2 _34462_ (.A(_05898_),
    .B(_05900_),
    .C(_06343_),
    .X(_06346_));
 sky130_fd_sc_hd__and2_2 _34463_ (.A(_06345_),
    .B(_06346_),
    .X(_06348_));
 sky130_fd_sc_hd__o21ai_2 _34464_ (.A1(_05859_),
    .A2(_05863_),
    .B1(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__or3_2 _34465_ (.A(_05859_),
    .B(_05863_),
    .C(_06348_),
    .X(_06350_));
 sky130_fd_sc_hd__nand2_2 _34466_ (.A(_06349_),
    .B(_06350_),
    .Y(_06351_));
 sky130_fd_sc_hd__o21bai_2 _34467_ (.A1(_05903_),
    .A2(_05905_),
    .B1_N(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__or3b_2 _34468_ (.A(_05903_),
    .B(_05905_),
    .C_N(_06351_),
    .X(_06353_));
 sky130_fd_sc_hd__nand2_2 _34469_ (.A(_06352_),
    .B(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__nand2_2 _34470_ (.A(_05907_),
    .B(_05909_),
    .Y(_06355_));
 sky130_fd_sc_hd__o21a_2 _34471_ (.A1(_05910_),
    .A2(_05911_),
    .B1(_06355_),
    .X(_06356_));
 sky130_fd_sc_hd__xor2_2 _34472_ (.A(_06354_),
    .B(_06356_),
    .X(_06357_));
 sky130_fd_sc_hd__xor2_2 _34473_ (.A(_06227_),
    .B(_06357_),
    .X(_06359_));
 sky130_fd_sc_hd__xnor2_2 _34474_ (.A(_06082_),
    .B(_06359_),
    .Y(_06360_));
 sky130_fd_sc_hd__a21oi_2 _34475_ (.A1(_06080_),
    .A2(_06081_),
    .B1(_06360_),
    .Y(_06361_));
 sky130_fd_sc_hd__and3_2 _34476_ (.A(_06080_),
    .B(_06081_),
    .C(_06360_),
    .X(_06362_));
 sky130_fd_sc_hd__nor2_2 _34477_ (.A(_06361_),
    .B(_06362_),
    .Y(_06363_));
 sky130_fd_sc_hd__and2_2 _34478_ (.A(_05758_),
    .B(_06067_),
    .X(_06364_));
 sky130_fd_sc_hd__inv_2 _34479_ (.A(_06364_),
    .Y(_06365_));
 sky130_fd_sc_hd__nor2_2 _34480_ (.A(_06065_),
    .B(_06066_),
    .Y(_06366_));
 sky130_fd_sc_hd__nand2_2 _34481_ (.A(_06065_),
    .B(_06066_),
    .Y(_06367_));
 sky130_fd_sc_hd__o21a_2 _34482_ (.A1(_06068_),
    .A2(_06366_),
    .B1(_06367_),
    .X(_06368_));
 sky130_fd_sc_hd__o21ba_2 _34483_ (.A1(_05767_),
    .A2(_06365_),
    .B1_N(_06368_),
    .X(_06370_));
 sky130_fd_sc_hd__xnor2_2 _34484_ (.A(_06363_),
    .B(_06370_),
    .Y(_06371_));
 sky130_fd_sc_hd__xnor2_2 _34485_ (.A(_13831_),
    .B(_06371_),
    .Y(_06372_));
 sky130_fd_sc_hd__and2b_2 _34486_ (.A_N(_06079_),
    .B(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__and2b_2 _34487_ (.A_N(_06372_),
    .B(_06079_),
    .X(_06374_));
 sky130_fd_sc_hd__nor2_2 _34488_ (.A(_06373_),
    .B(_06374_),
    .Y(oO[74]));
 sky130_fd_sc_hd__inv_2 _34489_ (.A(_06363_),
    .Y(_06375_));
 sky130_fd_sc_hd__o21ba_2 _34490_ (.A1(_06375_),
    .A2(_06370_),
    .B1_N(_06361_),
    .X(_06376_));
 sky130_fd_sc_hd__nor2_2 _34491_ (.A(_06227_),
    .B(_06357_),
    .Y(_06377_));
 sky130_fd_sc_hd__a21o_2 _34492_ (.A1(_06082_),
    .A2(_06359_),
    .B1(_06377_),
    .X(_06378_));
 sky130_fd_sc_hd__or2_2 _34493_ (.A(_06219_),
    .B(_06220_),
    .X(_06380_));
 sky130_fd_sc_hd__o21ai_2 _34494_ (.A1(_06221_),
    .A2(_06225_),
    .B1(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__or2b_2 _34495_ (.A(_06214_),
    .B_N(_06217_),
    .X(_06382_));
 sky130_fd_sc_hd__nand2_2 _34496_ (.A(_05920_),
    .B(_06218_),
    .Y(_06383_));
 sky130_fd_sc_hd__or2b_2 _34497_ (.A(_06209_),
    .B_N(_06212_),
    .X(_06384_));
 sky130_fd_sc_hd__nand2_2 _34498_ (.A(_06091_),
    .B(_06213_),
    .Y(_06385_));
 sky130_fd_sc_hd__and2_2 _34499_ (.A(_06205_),
    .B(_06207_),
    .X(_06386_));
 sky130_fd_sc_hd__nor2_2 _34500_ (.A(_06142_),
    .B(_06208_),
    .Y(_06387_));
 sky130_fd_sc_hd__nand2_2 _34501_ (.A(_06143_),
    .B(_06161_),
    .Y(_06388_));
 sky130_fd_sc_hd__or2_2 _34502_ (.A(_06162_),
    .B(_06203_),
    .X(_06389_));
 sky130_fd_sc_hd__and2_2 _34503_ (.A(_06148_),
    .B(_06159_),
    .X(_06391_));
 sky130_fd_sc_hd__a22o_2 _34504_ (.A1(_03023_),
    .A2(_03458_),
    .B1(_04905_),
    .B2(_14593_),
    .X(_06392_));
 sky130_fd_sc_hd__or3_2 _34505_ (.A(_01028_),
    .B(_05550_),
    .C(_06150_),
    .X(_06393_));
 sky130_fd_sc_hd__and2_2 _34506_ (.A(_06392_),
    .B(_06393_),
    .X(_06394_));
 sky130_fd_sc_hd__nor2_2 _34507_ (.A(_17672_),
    .B(_03068_),
    .Y(_06395_));
 sky130_fd_sc_hd__o22a_2 _34508_ (.A1(_01576_),
    .A2(_04181_),
    .B1(_04901_),
    .B2(_02608_),
    .X(_06396_));
 sky130_fd_sc_hd__or2_2 _34509_ (.A(_06395_),
    .B(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__a211o_2 _34510_ (.A1(_05209_),
    .A2(_05215_),
    .B1(_06038_),
    .C1(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__buf_1 _34511_ (.A(_03068_),
    .X(_06399_));
 sky130_fd_sc_hd__o22a_2 _34512_ (.A1(_16647_),
    .A2(_06399_),
    .B1(_06144_),
    .B2(_06146_),
    .X(_06400_));
 sky130_fd_sc_hd__o22ai_2 _34513_ (.A1(_06145_),
    .A2(_06398_),
    .B1(_06400_),
    .B2(_06397_),
    .Y(_06402_));
 sky130_fd_sc_hd__inv_2 _34514_ (.A(_06402_),
    .Y(_06403_));
 sky130_fd_sc_hd__o221ai_2 _34515_ (.A1(_16647_),
    .A2(_06399_),
    .B1(_06145_),
    .B2(_06147_),
    .C1(_06397_),
    .Y(_06404_));
 sky130_fd_sc_hd__nand3_2 _34516_ (.A(_06394_),
    .B(_06403_),
    .C(_06404_),
    .Y(_06405_));
 sky130_fd_sc_hd__a21o_2 _34517_ (.A1(_06403_),
    .A2(_06404_),
    .B1(_06394_),
    .X(_06406_));
 sky130_fd_sc_hd__and3_2 _34518_ (.A(_06391_),
    .B(_06405_),
    .C(_06406_),
    .X(_06407_));
 sky130_fd_sc_hd__a21oi_2 _34519_ (.A1(_06405_),
    .A2(_06406_),
    .B1(_06391_),
    .Y(_06408_));
 sky130_fd_sc_hd__a21o_2 _34520_ (.A1(_06181_),
    .A2(_06198_),
    .B1(_06196_),
    .X(_06409_));
 sky130_fd_sc_hd__or3_2 _34521_ (.A(_05978_),
    .B(_05504_),
    .C(_06165_),
    .X(_06410_));
 sky130_fd_sc_hd__buf_1 _34522_ (.A(_02984_),
    .X(_06411_));
 sky130_fd_sc_hd__buf_1 _34523_ (.A(_00662_),
    .X(_06413_));
 sky130_fd_sc_hd__buf_1 _34524_ (.A(_17394_),
    .X(_06414_));
 sky130_fd_sc_hd__a22o_2 _34525_ (.A1(_06411_),
    .A2(_03973_),
    .B1(_06413_),
    .B2(_06414_),
    .X(_06415_));
 sky130_fd_sc_hd__and2_2 _34526_ (.A(_06410_),
    .B(_06415_),
    .X(_06416_));
 sky130_fd_sc_hd__nor2_2 _34527_ (.A(_05979_),
    .B(_05500_),
    .Y(_06417_));
 sky130_fd_sc_hd__xnor2_2 _34528_ (.A(_06416_),
    .B(_06417_),
    .Y(_06418_));
 sky130_fd_sc_hd__nor2_2 _34529_ (.A(_16258_),
    .B(_01070_),
    .Y(_06419_));
 sky130_fd_sc_hd__o22a_2 _34530_ (.A1(_16606_),
    .A2(_04162_),
    .B1(_01070_),
    .B2(_01804_),
    .X(_06420_));
 sky130_fd_sc_hd__a21oi_2 _34531_ (.A1(_06169_),
    .A2(_06419_),
    .B1(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__nor2_2 _34532_ (.A(_04847_),
    .B(_05522_),
    .Y(_06422_));
 sky130_fd_sc_hd__xnor2_2 _34533_ (.A(_06421_),
    .B(_06422_),
    .Y(_06424_));
 sky130_fd_sc_hd__a21bo_2 _34534_ (.A1(_06173_),
    .A2(_06174_),
    .B1_N(_06170_),
    .X(_06425_));
 sky130_fd_sc_hd__or2b_2 _34535_ (.A(_06424_),
    .B_N(_06425_),
    .X(_06426_));
 sky130_fd_sc_hd__or2b_2 _34536_ (.A(_06425_),
    .B_N(_06424_),
    .X(_06427_));
 sky130_fd_sc_hd__nand2_2 _34537_ (.A(_06426_),
    .B(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__xnor2_2 _34538_ (.A(_06418_),
    .B(_06428_),
    .Y(_06429_));
 sky130_fd_sc_hd__a21o_2 _34539_ (.A1(_06188_),
    .A2(_06189_),
    .B1(_06186_),
    .X(_06430_));
 sky130_fd_sc_hd__and3_2 _34540_ (.A(_14593_),
    .B(_03458_),
    .C(_06151_),
    .X(_06431_));
 sky130_fd_sc_hd__nor2_2 _34541_ (.A(_14949_),
    .B(_02391_),
    .Y(_06432_));
 sky130_fd_sc_hd__xor2_2 _34542_ (.A(_06185_),
    .B(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__and3b_2 _34543_ (.A_N(_05521_),
    .B(_03438_),
    .C(_06433_),
    .X(_06435_));
 sky130_fd_sc_hd__o21ba_2 _34544_ (.A1(_05521_),
    .A2(_05543_),
    .B1_N(_06433_),
    .X(_06436_));
 sky130_fd_sc_hd__nor2_2 _34545_ (.A(_06435_),
    .B(_06436_),
    .Y(_06437_));
 sky130_fd_sc_hd__o21a_2 _34546_ (.A1(_06431_),
    .A2(_06153_),
    .B1(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__nor3_2 _34547_ (.A(_06431_),
    .B(_06153_),
    .C(_06437_),
    .Y(_06439_));
 sky130_fd_sc_hd__nor2_2 _34548_ (.A(_06438_),
    .B(_06439_),
    .Y(_06440_));
 sky130_fd_sc_hd__xnor2_2 _34549_ (.A(_06430_),
    .B(_06440_),
    .Y(_06441_));
 sky130_fd_sc_hd__a21bo_2 _34550_ (.A1(_06184_),
    .A2(_06192_),
    .B1_N(_06191_),
    .X(_06442_));
 sky130_fd_sc_hd__xor2_2 _34551_ (.A(_06441_),
    .B(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__xnor2_2 _34552_ (.A(_06429_),
    .B(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__nor2_2 _34553_ (.A(_06157_),
    .B(_06444_),
    .Y(_06446_));
 sky130_fd_sc_hd__and2_2 _34554_ (.A(_06157_),
    .B(_06444_),
    .X(_06447_));
 sky130_fd_sc_hd__nor2_2 _34555_ (.A(_06446_),
    .B(_06447_),
    .Y(_06448_));
 sky130_fd_sc_hd__xor2_2 _34556_ (.A(_06409_),
    .B(_06448_),
    .X(_06449_));
 sky130_fd_sc_hd__nor3b_2 _34557_ (.A(_06407_),
    .B(_06408_),
    .C_N(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__o21ba_2 _34558_ (.A1(_06407_),
    .A2(_06408_),
    .B1_N(_06449_),
    .X(_06451_));
 sky130_fd_sc_hd__a211oi_2 _34559_ (.A1(_06388_),
    .A2(_06389_),
    .B1(_06450_),
    .C1(_06451_),
    .Y(_06452_));
 sky130_fd_sc_hd__o211a_2 _34560_ (.A1(_06450_),
    .A2(_06451_),
    .B1(_06388_),
    .C1(_06389_),
    .X(_06453_));
 sky130_fd_sc_hd__o21ai_2 _34561_ (.A1(_06135_),
    .A2(_06136_),
    .B1(_06134_),
    .Y(_06454_));
 sky130_fd_sc_hd__or2b_2 _34562_ (.A(_06119_),
    .B_N(_06139_),
    .X(_06455_));
 sky130_fd_sc_hd__nand2_2 _34563_ (.A(_06454_),
    .B(_06455_),
    .Y(_06457_));
 sky130_fd_sc_hd__a21o_2 _34564_ (.A1(_06164_),
    .A2(_06202_),
    .B1(_06200_),
    .X(_06458_));
 sky130_fd_sc_hd__o31ai_2 _34565_ (.A1(_01576_),
    .A2(_05441_),
    .A3(_06099_),
    .B1(_06097_),
    .Y(_06459_));
 sky130_fd_sc_hd__nand2_2 _34566_ (.A(_02994_),
    .B(_02928_),
    .Y(_06460_));
 sky130_fd_sc_hd__or3_2 _34567_ (.A(_02463_),
    .B(_02317_),
    .C(_06460_),
    .X(_06461_));
 sky130_fd_sc_hd__o21ai_2 _34568_ (.A1(_02463_),
    .A2(_02317_),
    .B1(_06460_),
    .Y(_06462_));
 sky130_fd_sc_hd__nand2_2 _34569_ (.A(_06461_),
    .B(_06462_),
    .Y(_06463_));
 sky130_fd_sc_hd__nor2_2 _34570_ (.A(_01583_),
    .B(_03318_),
    .Y(_06464_));
 sky130_fd_sc_hd__xnor2_2 _34571_ (.A(_06463_),
    .B(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__nand2_2 _34572_ (.A(_01040_),
    .B(_01757_),
    .Y(_06466_));
 sky130_fd_sc_hd__xnor2_2 _34573_ (.A(_06102_),
    .B(_06466_),
    .Y(_06468_));
 sky130_fd_sc_hd__nand2_2 _34574_ (.A(_02989_),
    .B(_03327_),
    .Y(_06469_));
 sky130_fd_sc_hd__xnor2_2 _34575_ (.A(_06468_),
    .B(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__o22a_2 _34576_ (.A1(_05936_),
    .A2(_06102_),
    .B1(_06103_),
    .B2(_06106_),
    .X(_06471_));
 sky130_fd_sc_hd__nor2_2 _34577_ (.A(_06470_),
    .B(_06471_),
    .Y(_06472_));
 sky130_fd_sc_hd__nand2_2 _34578_ (.A(_06470_),
    .B(_06471_),
    .Y(_06473_));
 sky130_fd_sc_hd__and2b_2 _34579_ (.A_N(_06472_),
    .B(_06473_),
    .X(_06474_));
 sky130_fd_sc_hd__xnor2_2 _34580_ (.A(_06465_),
    .B(_06474_),
    .Y(_06475_));
 sky130_fd_sc_hd__a21oi_2 _34581_ (.A1(_06110_),
    .A2(_06113_),
    .B1(_06475_),
    .Y(_06476_));
 sky130_fd_sc_hd__and3_2 _34582_ (.A(_06110_),
    .B(_06113_),
    .C(_06475_),
    .X(_06477_));
 sky130_fd_sc_hd__nor2_2 _34583_ (.A(_06476_),
    .B(_06477_),
    .Y(_06479_));
 sky130_fd_sc_hd__xnor2_2 _34584_ (.A(_06459_),
    .B(_06479_),
    .Y(_06480_));
 sky130_fd_sc_hd__or2b_2 _34585_ (.A(_06130_),
    .B_N(_06124_),
    .X(_06481_));
 sky130_fd_sc_hd__a21bo_2 _34586_ (.A1(_06123_),
    .A2(_06131_),
    .B1_N(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__o21a_2 _34587_ (.A1(_06168_),
    .A2(_06180_),
    .B1(_06178_),
    .X(_06483_));
 sky130_fd_sc_hd__buf_1 _34588_ (.A(_04469_),
    .X(_06484_));
 sky130_fd_sc_hd__a31o_2 _34589_ (.A1(_01040_),
    .A2(_06484_),
    .A3(_06128_),
    .B1(_06125_),
    .X(_06485_));
 sky130_fd_sc_hd__nor2_2 _34590_ (.A(_05976_),
    .B(_06165_),
    .Y(_06486_));
 sky130_fd_sc_hd__a31o_2 _34591_ (.A1(_03024_),
    .A2(_03345_),
    .A3(_06166_),
    .B1(_06486_),
    .X(_06487_));
 sky130_fd_sc_hd__buf_1 _34592_ (.A(_18734_),
    .X(_06488_));
 sky130_fd_sc_hd__and4_2 _34593_ (.A(_01837_),
    .B(_03024_),
    .C(_18328_),
    .D(_06488_),
    .X(_06490_));
 sky130_fd_sc_hd__buf_1 _34594_ (.A(_18114_),
    .X(_06491_));
 sky130_fd_sc_hd__o22a_2 _34595_ (.A1(_04501_),
    .A2(_06491_),
    .B1(_18343_),
    .B2(_05983_),
    .X(_06492_));
 sky130_fd_sc_hd__nor2_2 _34596_ (.A(_06490_),
    .B(_06492_),
    .Y(_06493_));
 sky130_fd_sc_hd__nand2_2 _34597_ (.A(_04837_),
    .B(_04469_),
    .Y(_06494_));
 sky130_fd_sc_hd__xor2_2 _34598_ (.A(_06493_),
    .B(_06494_),
    .X(_06495_));
 sky130_fd_sc_hd__xnor2_2 _34599_ (.A(_06487_),
    .B(_06495_),
    .Y(_06496_));
 sky130_fd_sc_hd__xnor2_2 _34600_ (.A(_06485_),
    .B(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__xnor2_2 _34601_ (.A(_06483_),
    .B(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__xnor2_2 _34602_ (.A(_06482_),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__nor2_2 _34603_ (.A(_06122_),
    .B(_06132_),
    .Y(_06501_));
 sky130_fd_sc_hd__and2b_2 _34604_ (.A_N(_06133_),
    .B(_06121_),
    .X(_06502_));
 sky130_fd_sc_hd__nor2_2 _34605_ (.A(_06501_),
    .B(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__xnor2_2 _34606_ (.A(_06499_),
    .B(_06503_),
    .Y(_06504_));
 sky130_fd_sc_hd__xnor2_2 _34607_ (.A(_06480_),
    .B(_06504_),
    .Y(_06505_));
 sky130_fd_sc_hd__xnor2_2 _34608_ (.A(_06458_),
    .B(_06505_),
    .Y(_06506_));
 sky130_fd_sc_hd__xor2_2 _34609_ (.A(_06457_),
    .B(_06506_),
    .X(_06507_));
 sky130_fd_sc_hd__or3_2 _34610_ (.A(_06452_),
    .B(_06453_),
    .C(_06507_),
    .X(_06508_));
 sky130_fd_sc_hd__o21ai_2 _34611_ (.A1(_06452_),
    .A2(_06453_),
    .B1(_06507_),
    .Y(_06509_));
 sky130_fd_sc_hd__o211a_2 _34612_ (.A1(_06386_),
    .A2(_06387_),
    .B1(_06508_),
    .C1(_06509_),
    .X(_06510_));
 sky130_fd_sc_hd__a211oi_2 _34613_ (.A1(_06508_),
    .A2(_06509_),
    .B1(_06386_),
    .C1(_06387_),
    .Y(_06512_));
 sky130_fd_sc_hd__nand2_2 _34614_ (.A(_06095_),
    .B(_06140_),
    .Y(_06513_));
 sky130_fd_sc_hd__or2b_2 _34615_ (.A(_06141_),
    .B_N(_06093_),
    .X(_06514_));
 sky130_fd_sc_hd__a32oi_2 _34616_ (.A1(_06113_),
    .A2(_06114_),
    .A3(_06117_),
    .B1(_06118_),
    .B2(_06096_),
    .Y(_06515_));
 sky130_fd_sc_hd__a21oi_2 _34617_ (.A1(_06513_),
    .A2(_06514_),
    .B1(_06515_),
    .Y(_06516_));
 sky130_fd_sc_hd__and3_2 _34618_ (.A(_06513_),
    .B(_06514_),
    .C(_06515_),
    .X(_06517_));
 sky130_fd_sc_hd__nor2_2 _34619_ (.A(_06516_),
    .B(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__nor3b_2 _34620_ (.A(_06510_),
    .B(_06512_),
    .C_N(_06518_),
    .Y(_06519_));
 sky130_fd_sc_hd__o21ba_2 _34621_ (.A1(_06510_),
    .A2(_06512_),
    .B1_N(_06518_),
    .X(_06520_));
 sky130_fd_sc_hd__a211o_2 _34622_ (.A1(_06384_),
    .A2(_06385_),
    .B1(_06519_),
    .C1(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__o211ai_2 _34623_ (.A1(_06519_),
    .A2(_06520_),
    .B1(_06384_),
    .C1(_06385_),
    .Y(_06523_));
 sky130_fd_sc_hd__and3_2 _34624_ (.A(_06089_),
    .B(_06521_),
    .C(_06523_),
    .X(_06524_));
 sky130_fd_sc_hd__a21oi_2 _34625_ (.A1(_06521_),
    .A2(_06523_),
    .B1(_06089_),
    .Y(_06525_));
 sky130_fd_sc_hd__a211oi_2 _34626_ (.A1(_06382_),
    .A2(_06383_),
    .B1(_06524_),
    .C1(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__o211a_2 _34627_ (.A1(_06524_),
    .A2(_06525_),
    .B1(_06382_),
    .C1(_06383_),
    .X(_06527_));
 sky130_fd_sc_hd__nor2_2 _34628_ (.A(_06526_),
    .B(_06527_),
    .Y(_06528_));
 sky130_fd_sc_hd__xnor2_2 _34629_ (.A(_06381_),
    .B(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__a21oi_2 _34630_ (.A1(_06228_),
    .A2(_06235_),
    .B1(_05784_),
    .Y(_06530_));
 sky130_fd_sc_hd__and3_2 _34631_ (.A(iY[44]),
    .B(iX[63]),
    .C(_06229_),
    .X(_06531_));
 sky130_fd_sc_hd__a21oi_2 _34632_ (.A1(iY[44]),
    .A2(iX[63]),
    .B1(_06229_),
    .Y(_06532_));
 sky130_fd_sc_hd__o2bb2a_2 _34633_ (.A1_N(iY[46]),
    .A2_N(iX[61]),
    .B1(_06531_),
    .B2(_06532_),
    .X(_06534_));
 sky130_fd_sc_hd__and4bb_2 _34634_ (.A_N(_06531_),
    .B_N(_06532_),
    .C(iY[46]),
    .D(iX[61]),
    .X(_06535_));
 sky130_fd_sc_hd__nor2_2 _34635_ (.A(_06534_),
    .B(_06535_),
    .Y(_06536_));
 sky130_fd_sc_hd__and2b_2 _34636_ (.A_N(_06530_),
    .B(_06536_),
    .X(_06537_));
 sky130_fd_sc_hd__and2b_2 _34637_ (.A_N(_06536_),
    .B(_06530_),
    .X(_06538_));
 sky130_fd_sc_hd__nor2_2 _34638_ (.A(_06537_),
    .B(_06538_),
    .Y(_06539_));
 sky130_fd_sc_hd__a21o_2 _34639_ (.A1(_05827_),
    .A2(_06258_),
    .B1(_06269_),
    .X(_06540_));
 sky130_fd_sc_hd__and2b_2 _34640_ (.A_N(_06236_),
    .B(_06239_),
    .X(_06541_));
 sky130_fd_sc_hd__and4_2 _34641_ (.A(iX[53]),
    .B(iY[53]),
    .C(iX[54]),
    .D(iY[54]),
    .X(_06542_));
 sky130_fd_sc_hd__a22oi_2 _34642_ (.A1(iY[53]),
    .A2(iX[54]),
    .B1(iY[54]),
    .B2(iX[53]),
    .Y(_06543_));
 sky130_fd_sc_hd__nor2_2 _34643_ (.A(_06542_),
    .B(_06543_),
    .Y(_06545_));
 sky130_fd_sc_hd__nand2_2 _34644_ (.A(iX[52]),
    .B(iY[55]),
    .Y(_06546_));
 sky130_fd_sc_hd__xnor2_2 _34645_ (.A(_06545_),
    .B(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__and4_2 _34646_ (.A(iY[50]),
    .B(iY[51]),
    .C(iX[56]),
    .D(iX[57]),
    .X(_06548_));
 sky130_fd_sc_hd__a22oi_2 _34647_ (.A1(iY[51]),
    .A2(iX[56]),
    .B1(iX[57]),
    .B2(iY[50]),
    .Y(_06549_));
 sky130_fd_sc_hd__nor2_2 _34648_ (.A(_06548_),
    .B(_06549_),
    .Y(_06550_));
 sky130_fd_sc_hd__nand2_2 _34649_ (.A(iY[52]),
    .B(iX[55]),
    .Y(_06551_));
 sky130_fd_sc_hd__xnor2_2 _34650_ (.A(_06550_),
    .B(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__o21ba_2 _34651_ (.A1(_06249_),
    .A2(_06251_),
    .B1_N(_06247_),
    .X(_06553_));
 sky130_fd_sc_hd__xnor2_2 _34652_ (.A(_06552_),
    .B(_06553_),
    .Y(_06554_));
 sky130_fd_sc_hd__and2_2 _34653_ (.A(_06547_),
    .B(_06554_),
    .X(_06556_));
 sky130_fd_sc_hd__nor2_2 _34654_ (.A(_06547_),
    .B(_06554_),
    .Y(_06557_));
 sky130_fd_sc_hd__or2_2 _34655_ (.A(_06556_),
    .B(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__or2b_2 _34656_ (.A(_06260_),
    .B_N(_06265_),
    .X(_06559_));
 sky130_fd_sc_hd__a31o_2 _34657_ (.A1(iY[49]),
    .A2(iX[57]),
    .A3(_06263_),
    .B1(_06261_),
    .X(_06560_));
 sky130_fd_sc_hd__and4_2 _34658_ (.A(iY[47]),
    .B(iY[48]),
    .C(iX[59]),
    .D(iX[60]),
    .X(_06561_));
 sky130_fd_sc_hd__a22oi_2 _34659_ (.A1(iY[48]),
    .A2(iX[59]),
    .B1(iX[60]),
    .B2(iY[47]),
    .Y(_06562_));
 sky130_fd_sc_hd__nor2_2 _34660_ (.A(_06561_),
    .B(_06562_),
    .Y(_06563_));
 sky130_fd_sc_hd__nand2_2 _34661_ (.A(iY[49]),
    .B(iX[58]),
    .Y(_06564_));
 sky130_fd_sc_hd__xnor2_2 _34662_ (.A(_06563_),
    .B(_06564_),
    .Y(_06565_));
 sky130_fd_sc_hd__o21ai_2 _34663_ (.A1(_06230_),
    .A2(_06234_),
    .B1(_06565_),
    .Y(_06567_));
 sky130_fd_sc_hd__or3_2 _34664_ (.A(_06230_),
    .B(_06234_),
    .C(_06565_),
    .X(_06568_));
 sky130_fd_sc_hd__and2_2 _34665_ (.A(_06567_),
    .B(_06568_),
    .X(_06569_));
 sky130_fd_sc_hd__xnor2_2 _34666_ (.A(_06560_),
    .B(_06569_),
    .Y(_06570_));
 sky130_fd_sc_hd__a21oi_2 _34667_ (.A1(_06559_),
    .A2(_06267_),
    .B1(_06570_),
    .Y(_06571_));
 sky130_fd_sc_hd__and3_2 _34668_ (.A(_06559_),
    .B(_06267_),
    .C(_06570_),
    .X(_06572_));
 sky130_fd_sc_hd__or3_2 _34669_ (.A(_06558_),
    .B(_06571_),
    .C(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__o21ai_2 _34670_ (.A1(_06571_),
    .A2(_06572_),
    .B1(_06558_),
    .Y(_06574_));
 sky130_fd_sc_hd__and3_2 _34671_ (.A(_06541_),
    .B(_06573_),
    .C(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__a21oi_2 _34672_ (.A1(_06573_),
    .A2(_06574_),
    .B1(_06541_),
    .Y(_06576_));
 sky130_fd_sc_hd__a211o_2 _34673_ (.A1(_06540_),
    .A2(_06273_),
    .B1(_06575_),
    .C1(_06576_),
    .X(_06578_));
 sky130_fd_sc_hd__o211ai_2 _34674_ (.A1(_06575_),
    .A2(_06576_),
    .B1(_06540_),
    .C1(_06273_),
    .Y(_06579_));
 sky130_fd_sc_hd__and3_2 _34675_ (.A(_06539_),
    .B(_06578_),
    .C(_06579_),
    .X(_06580_));
 sky130_fd_sc_hd__a21oi_2 _34676_ (.A1(_06578_),
    .A2(_06579_),
    .B1(_06539_),
    .Y(_06581_));
 sky130_fd_sc_hd__o21ai_2 _34677_ (.A1(_06580_),
    .A2(_06581_),
    .B1(_06279_),
    .Y(_06582_));
 sky130_fd_sc_hd__or3_2 _34678_ (.A(_06279_),
    .B(_06580_),
    .C(_06581_),
    .X(_06583_));
 sky130_fd_sc_hd__inv_2 _34679_ (.A(_06326_),
    .Y(_06584_));
 sky130_fd_sc_hd__or2b_2 _34680_ (.A(_06291_),
    .B_N(_06290_),
    .X(_06585_));
 sky130_fd_sc_hd__and4_2 _34681_ (.A(iX[47]),
    .B(iX[48]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_06586_));
 sky130_fd_sc_hd__a22oi_2 _34682_ (.A1(iX[48]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[47]),
    .Y(_06587_));
 sky130_fd_sc_hd__nor2_2 _34683_ (.A(_06586_),
    .B(_06587_),
    .Y(_06589_));
 sky130_fd_sc_hd__nand2_2 _34684_ (.A(iX[46]),
    .B(iY[61]),
    .Y(_06590_));
 sky130_fd_sc_hd__xnor2_2 _34685_ (.A(_06589_),
    .B(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__o21ba_2 _34686_ (.A1(_06287_),
    .A2(_06289_),
    .B1_N(_06286_),
    .X(_06592_));
 sky130_fd_sc_hd__xnor2_2 _34687_ (.A(_06591_),
    .B(_06592_),
    .Y(_06593_));
 sky130_fd_sc_hd__and2_2 _34688_ (.A(iX[45]),
    .B(iY[62]),
    .X(_06594_));
 sky130_fd_sc_hd__or2_2 _34689_ (.A(_06593_),
    .B(_06594_),
    .X(_06595_));
 sky130_fd_sc_hd__nand2_2 _34690_ (.A(_06593_),
    .B(_06594_),
    .Y(_06596_));
 sky130_fd_sc_hd__nand2_2 _34691_ (.A(_06595_),
    .B(_06596_),
    .Y(_06597_));
 sky130_fd_sc_hd__a21oi_2 _34692_ (.A1(_06585_),
    .A2(_06296_),
    .B1(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__and3_2 _34693_ (.A(_06585_),
    .B(_06296_),
    .C(_06597_),
    .X(_06600_));
 sky130_fd_sc_hd__nor2_2 _34694_ (.A(_06598_),
    .B(_06600_),
    .Y(_06601_));
 sky130_fd_sc_hd__nand2_2 _34695_ (.A(iX[44]),
    .B(iY[63]),
    .Y(_06602_));
 sky130_fd_sc_hd__xnor2_2 _34696_ (.A(_06601_),
    .B(_06602_),
    .Y(_06603_));
 sky130_fd_sc_hd__or2b_2 _34697_ (.A(_06311_),
    .B_N(_06317_),
    .X(_06604_));
 sky130_fd_sc_hd__or2b_2 _34698_ (.A(_06310_),
    .B_N(_06318_),
    .X(_06605_));
 sky130_fd_sc_hd__and2b_2 _34699_ (.A_N(_06253_),
    .B(_06252_),
    .X(_06606_));
 sky130_fd_sc_hd__o21ba_2 _34700_ (.A1(_06313_),
    .A2(_06316_),
    .B1_N(_06312_),
    .X(_06607_));
 sky130_fd_sc_hd__o21ba_2 _34701_ (.A1(_06243_),
    .A2(_06245_),
    .B1_N(_06242_),
    .X(_06608_));
 sky130_fd_sc_hd__and4_2 _34702_ (.A(iX[50]),
    .B(iX[51]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_06609_));
 sky130_fd_sc_hd__a22oi_2 _34703_ (.A1(iX[51]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[50]),
    .Y(_06611_));
 sky130_fd_sc_hd__nor2_2 _34704_ (.A(_06609_),
    .B(_06611_),
    .Y(_06612_));
 sky130_fd_sc_hd__nand2_2 _34705_ (.A(iX[49]),
    .B(iY[58]),
    .Y(_06613_));
 sky130_fd_sc_hd__xnor2_2 _34706_ (.A(_06612_),
    .B(_06613_),
    .Y(_06614_));
 sky130_fd_sc_hd__xnor2_2 _34707_ (.A(_06608_),
    .B(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__xnor2_2 _34708_ (.A(_06607_),
    .B(_06615_),
    .Y(_06616_));
 sky130_fd_sc_hd__o21a_2 _34709_ (.A1(_06606_),
    .A2(_06255_),
    .B1(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__nor3_2 _34710_ (.A(_06606_),
    .B(_06255_),
    .C(_06616_),
    .Y(_06618_));
 sky130_fd_sc_hd__a211oi_2 _34711_ (.A1(_06604_),
    .A2(_06605_),
    .B1(_06617_),
    .C1(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__o211a_2 _34712_ (.A1(_06617_),
    .A2(_06618_),
    .B1(_06604_),
    .C1(_06605_),
    .X(_06620_));
 sky130_fd_sc_hd__nor2_2 _34713_ (.A(_06320_),
    .B(_06322_),
    .Y(_06622_));
 sky130_fd_sc_hd__or3_2 _34714_ (.A(_06619_),
    .B(_06620_),
    .C(_06622_),
    .X(_06623_));
 sky130_fd_sc_hd__o21ai_2 _34715_ (.A1(_06619_),
    .A2(_06620_),
    .B1(_06622_),
    .Y(_06624_));
 sky130_fd_sc_hd__and3_2 _34716_ (.A(_06603_),
    .B(_06623_),
    .C(_06624_),
    .X(_06625_));
 sky130_fd_sc_hd__a21oi_2 _34717_ (.A1(_06623_),
    .A2(_06624_),
    .B1(_06603_),
    .Y(_06626_));
 sky130_fd_sc_hd__nor2_2 _34718_ (.A(_06625_),
    .B(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__o21ai_2 _34719_ (.A1(_06275_),
    .A2(_06277_),
    .B1(_06627_),
    .Y(_06628_));
 sky130_fd_sc_hd__or3_2 _34720_ (.A(_06275_),
    .B(_06277_),
    .C(_06627_),
    .X(_06629_));
 sky130_fd_sc_hd__o211ai_2 _34721_ (.A1(_06584_),
    .A2(_06328_),
    .B1(_06628_),
    .C1(_06629_),
    .Y(_06630_));
 sky130_fd_sc_hd__a211o_2 _34722_ (.A1(_06628_),
    .A2(_06629_),
    .B1(_06584_),
    .C1(_06328_),
    .X(_06631_));
 sky130_fd_sc_hd__nand4_2 _34723_ (.A(_06582_),
    .B(_06583_),
    .C(_06630_),
    .D(_06631_),
    .Y(_06633_));
 sky130_fd_sc_hd__a22o_2 _34724_ (.A1(_06582_),
    .A2(_06583_),
    .B1(_06630_),
    .B2(_06631_),
    .X(_06634_));
 sky130_fd_sc_hd__nand2_2 _34725_ (.A(_06284_),
    .B(_06335_),
    .Y(_06635_));
 sky130_fd_sc_hd__and3_2 _34726_ (.A(_06633_),
    .B(_06634_),
    .C(_06635_),
    .X(_06636_));
 sky130_fd_sc_hd__a21oi_2 _34727_ (.A1(_06633_),
    .A2(_06634_),
    .B1(_06635_),
    .Y(_06637_));
 sky130_fd_sc_hd__a211oi_2 _34728_ (.A1(_06331_),
    .A2(_06333_),
    .B1(_06636_),
    .C1(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__o211a_2 _34729_ (.A1(_06636_),
    .A2(_06637_),
    .B1(_06331_),
    .C1(_06333_),
    .X(_06639_));
 sky130_fd_sc_hd__nor2_2 _34730_ (.A(_06638_),
    .B(_06639_),
    .Y(_06640_));
 sky130_fd_sc_hd__o21a_2 _34731_ (.A1(_06339_),
    .A2(_06341_),
    .B1(_06640_),
    .X(_06641_));
 sky130_fd_sc_hd__nor3_2 _34732_ (.A(_06339_),
    .B(_06341_),
    .C(_06640_),
    .Y(_06642_));
 sky130_fd_sc_hd__a211oi_2 _34733_ (.A1(_06299_),
    .A2(_06305_),
    .B1(_06641_),
    .C1(_06642_),
    .Y(_06644_));
 sky130_fd_sc_hd__o211a_2 _34734_ (.A1(_06641_),
    .A2(_06642_),
    .B1(_06299_),
    .C1(_06305_),
    .X(_06645_));
 sky130_fd_sc_hd__o211a_2 _34735_ (.A1(_06644_),
    .A2(_06645_),
    .B1(_06345_),
    .C1(_06349_),
    .X(_06646_));
 sky130_fd_sc_hd__a211oi_2 _34736_ (.A1(_06345_),
    .A2(_06349_),
    .B1(_06644_),
    .C1(_06645_),
    .Y(_06647_));
 sky130_fd_sc_hd__nor2_2 _34737_ (.A(_06646_),
    .B(_06647_),
    .Y(_06648_));
 sky130_fd_sc_hd__o21ai_2 _34738_ (.A1(_06354_),
    .A2(_06356_),
    .B1(_06352_),
    .Y(_06649_));
 sky130_fd_sc_hd__xnor2_2 _34739_ (.A(_06648_),
    .B(_06649_),
    .Y(_06650_));
 sky130_fd_sc_hd__xnor2_2 _34740_ (.A(_06529_),
    .B(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__xor2_2 _34741_ (.A(_14204_),
    .B(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__xor2_2 _34742_ (.A(_06378_),
    .B(_06652_),
    .X(_06653_));
 sky130_fd_sc_hd__xnor2_2 _34743_ (.A(_06376_),
    .B(_06653_),
    .Y(_06655_));
 sky130_fd_sc_hd__and2b_2 _34744_ (.A_N(_06655_),
    .B(_14070_),
    .X(_06656_));
 sky130_fd_sc_hd__and2b_2 _34745_ (.A_N(_14070_),
    .B(_06655_),
    .X(_06657_));
 sky130_fd_sc_hd__nor2_2 _34746_ (.A(_06656_),
    .B(_06657_),
    .Y(_06658_));
 sky130_fd_sc_hd__and2b_2 _34747_ (.A_N(_13831_),
    .B(_06371_),
    .X(_06659_));
 sky130_fd_sc_hd__nor2_2 _34748_ (.A(_06659_),
    .B(_06373_),
    .Y(_06660_));
 sky130_fd_sc_hd__xnor2_2 _34749_ (.A(_06658_),
    .B(_06660_),
    .Y(oO[75]));
 sky130_fd_sc_hd__a22oi_2 _34750_ (.A1(iY[46]),
    .A2(iX[62]),
    .B1(iX[63]),
    .B2(iY[45]),
    .Y(_06661_));
 sky130_fd_sc_hd__and3_2 _34751_ (.A(iY[46]),
    .B(iX[63]),
    .C(_06229_),
    .X(_06662_));
 sky130_fd_sc_hd__a21o_2 _34752_ (.A1(_06559_),
    .A2(_06267_),
    .B1(_06570_),
    .X(_06663_));
 sky130_fd_sc_hd__and4_2 _34753_ (.A(iY[53]),
    .B(iX[54]),
    .C(iY[54]),
    .D(iX[55]),
    .X(_06665_));
 sky130_fd_sc_hd__a22oi_2 _34754_ (.A1(iX[54]),
    .A2(iY[54]),
    .B1(iX[55]),
    .B2(iY[53]),
    .Y(_06666_));
 sky130_fd_sc_hd__nor2_2 _34755_ (.A(_06665_),
    .B(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__nand2_2 _34756_ (.A(iX[53]),
    .B(iY[55]),
    .Y(_06668_));
 sky130_fd_sc_hd__xnor2_2 _34757_ (.A(_06667_),
    .B(_06668_),
    .Y(_06669_));
 sky130_fd_sc_hd__and4_2 _34758_ (.A(iY[50]),
    .B(iY[51]),
    .C(iX[57]),
    .D(iX[58]),
    .X(_06670_));
 sky130_fd_sc_hd__a22oi_2 _34759_ (.A1(iY[51]),
    .A2(iX[57]),
    .B1(iX[58]),
    .B2(iY[50]),
    .Y(_06671_));
 sky130_fd_sc_hd__nor2_2 _34760_ (.A(_06670_),
    .B(_06671_),
    .Y(_06672_));
 sky130_fd_sc_hd__nand2_2 _34761_ (.A(iY[52]),
    .B(iX[56]),
    .Y(_06673_));
 sky130_fd_sc_hd__xnor2_2 _34762_ (.A(_06672_),
    .B(_06673_),
    .Y(_06674_));
 sky130_fd_sc_hd__o21ba_2 _34763_ (.A1(_06549_),
    .A2(_06551_),
    .B1_N(_06548_),
    .X(_06676_));
 sky130_fd_sc_hd__xnor2_2 _34764_ (.A(_06674_),
    .B(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__and2_2 _34765_ (.A(_06669_),
    .B(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__nor2_2 _34766_ (.A(_06669_),
    .B(_06677_),
    .Y(_06679_));
 sky130_fd_sc_hd__or2_2 _34767_ (.A(_06678_),
    .B(_06679_),
    .X(_06680_));
 sky130_fd_sc_hd__nand2_2 _34768_ (.A(_06560_),
    .B(_06569_),
    .Y(_06681_));
 sky130_fd_sc_hd__a31o_2 _34769_ (.A1(iY[49]),
    .A2(iX[58]),
    .A3(_06563_),
    .B1(_06561_),
    .X(_06682_));
 sky130_fd_sc_hd__and4_2 _34770_ (.A(iY[47]),
    .B(iY[48]),
    .C(iX[60]),
    .D(iX[61]),
    .X(_06683_));
 sky130_fd_sc_hd__a22oi_2 _34771_ (.A1(iY[48]),
    .A2(iX[60]),
    .B1(iX[61]),
    .B2(iY[47]),
    .Y(_06684_));
 sky130_fd_sc_hd__nor2_2 _34772_ (.A(_06683_),
    .B(_06684_),
    .Y(_06685_));
 sky130_fd_sc_hd__nand2_2 _34773_ (.A(iY[49]),
    .B(iX[59]),
    .Y(_06687_));
 sky130_fd_sc_hd__xnor2_2 _34774_ (.A(_06685_),
    .B(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__o21ai_2 _34775_ (.A1(_06531_),
    .A2(_06535_),
    .B1(_06688_),
    .Y(_06689_));
 sky130_fd_sc_hd__or3_2 _34776_ (.A(_06531_),
    .B(_06535_),
    .C(_06688_),
    .X(_06690_));
 sky130_fd_sc_hd__and2_2 _34777_ (.A(_06689_),
    .B(_06690_),
    .X(_06691_));
 sky130_fd_sc_hd__xnor2_2 _34778_ (.A(_06682_),
    .B(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__a21oi_2 _34779_ (.A1(_06567_),
    .A2(_06681_),
    .B1(_06692_),
    .Y(_06693_));
 sky130_fd_sc_hd__and3_2 _34780_ (.A(_06567_),
    .B(_06681_),
    .C(_06692_),
    .X(_06694_));
 sky130_fd_sc_hd__or3_2 _34781_ (.A(_06680_),
    .B(_06693_),
    .C(_06694_),
    .X(_06695_));
 sky130_fd_sc_hd__o21ai_2 _34782_ (.A1(_06693_),
    .A2(_06694_),
    .B1(_06680_),
    .Y(_06696_));
 sky130_fd_sc_hd__and3_2 _34783_ (.A(_06537_),
    .B(_06695_),
    .C(_06696_),
    .X(_06698_));
 sky130_fd_sc_hd__a21oi_2 _34784_ (.A1(_06695_),
    .A2(_06696_),
    .B1(_06537_),
    .Y(_06699_));
 sky130_fd_sc_hd__a211oi_2 _34785_ (.A1(_06663_),
    .A2(_06573_),
    .B1(_06698_),
    .C1(_06699_),
    .Y(_06700_));
 sky130_fd_sc_hd__o211a_2 _34786_ (.A1(_06698_),
    .A2(_06699_),
    .B1(_06663_),
    .C1(_06573_),
    .X(_06701_));
 sky130_fd_sc_hd__or4_2 _34787_ (.A(_06661_),
    .B(_06662_),
    .C(_06700_),
    .D(_06701_),
    .X(_06702_));
 sky130_fd_sc_hd__o22ai_2 _34788_ (.A1(_06661_),
    .A2(_06662_),
    .B1(_06700_),
    .B2(_06701_),
    .Y(_06703_));
 sky130_fd_sc_hd__a21o_2 _34789_ (.A1(_06702_),
    .A2(_06703_),
    .B1(_06580_),
    .X(_06704_));
 sky130_fd_sc_hd__nand3_2 _34790_ (.A(_06580_),
    .B(_06702_),
    .C(_06703_),
    .Y(_06705_));
 sky130_fd_sc_hd__inv_2 _34791_ (.A(_06625_),
    .Y(_06706_));
 sky130_fd_sc_hd__or2b_2 _34792_ (.A(_06575_),
    .B_N(_06578_),
    .X(_06707_));
 sky130_fd_sc_hd__and4_2 _34793_ (.A(iX[48]),
    .B(iX[49]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_06709_));
 sky130_fd_sc_hd__a22oi_2 _34794_ (.A1(iX[49]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[48]),
    .Y(_06710_));
 sky130_fd_sc_hd__nor2_2 _34795_ (.A(_06709_),
    .B(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__nand2_2 _34796_ (.A(iX[47]),
    .B(iY[61]),
    .Y(_06712_));
 sky130_fd_sc_hd__xnor2_2 _34797_ (.A(_06711_),
    .B(_06712_),
    .Y(_06713_));
 sky130_fd_sc_hd__o21ba_2 _34798_ (.A1(_06587_),
    .A2(_06590_),
    .B1_N(_06586_),
    .X(_06714_));
 sky130_fd_sc_hd__xnor2_2 _34799_ (.A(_06713_),
    .B(_06714_),
    .Y(_06715_));
 sky130_fd_sc_hd__and2_2 _34800_ (.A(iX[46]),
    .B(iY[62]),
    .X(_06716_));
 sky130_fd_sc_hd__or2_2 _34801_ (.A(_06715_),
    .B(_06716_),
    .X(_06717_));
 sky130_fd_sc_hd__nand2_2 _34802_ (.A(_06715_),
    .B(_06716_),
    .Y(_06718_));
 sky130_fd_sc_hd__nand2_2 _34803_ (.A(_06717_),
    .B(_06718_),
    .Y(_06720_));
 sky130_fd_sc_hd__or2b_2 _34804_ (.A(_06592_),
    .B_N(_06591_),
    .X(_06721_));
 sky130_fd_sc_hd__nand2_2 _34805_ (.A(_06721_),
    .B(_06596_),
    .Y(_06722_));
 sky130_fd_sc_hd__xnor2_2 _34806_ (.A(_06720_),
    .B(_06722_),
    .Y(_06723_));
 sky130_fd_sc_hd__and2_2 _34807_ (.A(iX[45]),
    .B(iY[63]),
    .X(_06724_));
 sky130_fd_sc_hd__nor2_2 _34808_ (.A(_06723_),
    .B(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__and2_2 _34809_ (.A(_06723_),
    .B(_06724_),
    .X(_06726_));
 sky130_fd_sc_hd__nor2_2 _34810_ (.A(_06725_),
    .B(_06726_),
    .Y(_06727_));
 sky130_fd_sc_hd__or2b_2 _34811_ (.A(_06608_),
    .B_N(_06614_),
    .X(_06728_));
 sky130_fd_sc_hd__or2b_2 _34812_ (.A(_06607_),
    .B_N(_06615_),
    .X(_06729_));
 sky130_fd_sc_hd__and2b_2 _34813_ (.A_N(_06553_),
    .B(_06552_),
    .X(_06731_));
 sky130_fd_sc_hd__o21ba_2 _34814_ (.A1(_06611_),
    .A2(_06613_),
    .B1_N(_06609_),
    .X(_06732_));
 sky130_fd_sc_hd__o21ba_2 _34815_ (.A1(_06543_),
    .A2(_06546_),
    .B1_N(_06542_),
    .X(_06733_));
 sky130_fd_sc_hd__and4_2 _34816_ (.A(iX[51]),
    .B(iX[52]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_06734_));
 sky130_fd_sc_hd__a22oi_2 _34817_ (.A1(iX[52]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[51]),
    .Y(_06735_));
 sky130_fd_sc_hd__nor2_2 _34818_ (.A(_06734_),
    .B(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__nand2_2 _34819_ (.A(iX[50]),
    .B(iY[58]),
    .Y(_06737_));
 sky130_fd_sc_hd__xnor2_2 _34820_ (.A(_06736_),
    .B(_06737_),
    .Y(_06738_));
 sky130_fd_sc_hd__xnor2_2 _34821_ (.A(_06733_),
    .B(_06738_),
    .Y(_06739_));
 sky130_fd_sc_hd__xnor2_2 _34822_ (.A(_06732_),
    .B(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__o21a_2 _34823_ (.A1(_06731_),
    .A2(_06556_),
    .B1(_06740_),
    .X(_06741_));
 sky130_fd_sc_hd__nor3_2 _34824_ (.A(_06731_),
    .B(_06556_),
    .C(_06740_),
    .Y(_06742_));
 sky130_fd_sc_hd__a211oi_2 _34825_ (.A1(_06728_),
    .A2(_06729_),
    .B1(_06741_),
    .C1(_06742_),
    .Y(_06743_));
 sky130_fd_sc_hd__o211a_2 _34826_ (.A1(_06741_),
    .A2(_06742_),
    .B1(_06728_),
    .C1(_06729_),
    .X(_06744_));
 sky130_fd_sc_hd__nor2_2 _34827_ (.A(_06617_),
    .B(_06619_),
    .Y(_06745_));
 sky130_fd_sc_hd__or3_2 _34828_ (.A(_06743_),
    .B(_06744_),
    .C(_06745_),
    .X(_06746_));
 sky130_fd_sc_hd__o21ai_2 _34829_ (.A1(_06743_),
    .A2(_06744_),
    .B1(_06745_),
    .Y(_06747_));
 sky130_fd_sc_hd__and3_2 _34830_ (.A(_06727_),
    .B(_06746_),
    .C(_06747_),
    .X(_06748_));
 sky130_fd_sc_hd__a21oi_2 _34831_ (.A1(_06746_),
    .A2(_06747_),
    .B1(_06727_),
    .Y(_06749_));
 sky130_fd_sc_hd__nor2_2 _34832_ (.A(_06748_),
    .B(_06749_),
    .Y(_06750_));
 sky130_fd_sc_hd__xnor2_2 _34833_ (.A(_06707_),
    .B(_06750_),
    .Y(_06752_));
 sky130_fd_sc_hd__a21o_2 _34834_ (.A1(_06623_),
    .A2(_06706_),
    .B1(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__nand3_2 _34835_ (.A(_06623_),
    .B(_06706_),
    .C(_06752_),
    .Y(_06754_));
 sky130_fd_sc_hd__nand4_2 _34836_ (.A(_06704_),
    .B(_06705_),
    .C(_06753_),
    .D(_06754_),
    .Y(_06755_));
 sky130_fd_sc_hd__a22o_2 _34837_ (.A1(_06704_),
    .A2(_06705_),
    .B1(_06753_),
    .B2(_06754_),
    .X(_06756_));
 sky130_fd_sc_hd__nand2_2 _34838_ (.A(_06583_),
    .B(_06633_),
    .Y(_06757_));
 sky130_fd_sc_hd__and3_2 _34839_ (.A(_06755_),
    .B(_06756_),
    .C(_06757_),
    .X(_06758_));
 sky130_fd_sc_hd__a21oi_2 _34840_ (.A1(_06755_),
    .A2(_06756_),
    .B1(_06757_),
    .Y(_06759_));
 sky130_fd_sc_hd__or2_2 _34841_ (.A(_06758_),
    .B(_06759_),
    .X(_06760_));
 sky130_fd_sc_hd__nand2_2 _34842_ (.A(_06628_),
    .B(_06630_),
    .Y(_06761_));
 sky130_fd_sc_hd__xnor2_2 _34843_ (.A(_06760_),
    .B(_06761_),
    .Y(_06763_));
 sky130_fd_sc_hd__nor2_2 _34844_ (.A(_06636_),
    .B(_06638_),
    .Y(_06764_));
 sky130_fd_sc_hd__xnor2_2 _34845_ (.A(_06763_),
    .B(_06764_),
    .Y(_06765_));
 sky130_fd_sc_hd__a31o_2 _34846_ (.A1(iX[44]),
    .A2(iY[63]),
    .A3(_06601_),
    .B1(_06598_),
    .X(_06766_));
 sky130_fd_sc_hd__xnor2_2 _34847_ (.A(_06765_),
    .B(_06766_),
    .Y(_06767_));
 sky130_fd_sc_hd__nor2_2 _34848_ (.A(_06641_),
    .B(_06644_),
    .Y(_06768_));
 sky130_fd_sc_hd__nor2_2 _34849_ (.A(_06767_),
    .B(_06768_),
    .Y(_06769_));
 sky130_fd_sc_hd__and2_2 _34850_ (.A(_06767_),
    .B(_06768_),
    .X(_06770_));
 sky130_fd_sc_hd__nor2_2 _34851_ (.A(_06769_),
    .B(_06770_),
    .Y(_06771_));
 sky130_fd_sc_hd__or3b_2 _34852_ (.A(_05910_),
    .B(_06354_),
    .C_N(_06648_),
    .X(_06772_));
 sky130_fd_sc_hd__a2111o_2 _34853_ (.A1(_05086_),
    .A2(_05594_),
    .B1(_05595_),
    .C1(_06772_),
    .D1(_05746_),
    .X(_06774_));
 sky130_fd_sc_hd__o21a_2 _34854_ (.A1(_05743_),
    .A2(_05910_),
    .B1(_06355_),
    .X(_06775_));
 sky130_fd_sc_hd__or3b_2 _34855_ (.A(_06354_),
    .B(_06775_),
    .C_N(_06648_),
    .X(_06776_));
 sky130_fd_sc_hd__or2_2 _34856_ (.A(_06352_),
    .B(_06646_),
    .X(_06777_));
 sky130_fd_sc_hd__and3b_2 _34857_ (.A_N(_06647_),
    .B(_06776_),
    .C(_06777_),
    .X(_06778_));
 sky130_fd_sc_hd__and2_2 _34858_ (.A(_06774_),
    .B(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__xnor2_2 _34859_ (.A(_06771_),
    .B(_06779_),
    .Y(_06780_));
 sky130_fd_sc_hd__nand3_2 _34860_ (.A(_06089_),
    .B(_06521_),
    .C(_06523_),
    .Y(_06781_));
 sky130_fd_sc_hd__nor3_2 _34861_ (.A(_06452_),
    .B(_06453_),
    .C(_06507_),
    .Y(_06782_));
 sky130_fd_sc_hd__buf_1 _34862_ (.A(_04905_),
    .X(_06783_));
 sky130_fd_sc_hd__or2_2 _34863_ (.A(_18405_),
    .B(_03068_),
    .X(_06785_));
 sky130_fd_sc_hd__buf_1 _34864_ (.A(_04181_),
    .X(_06786_));
 sky130_fd_sc_hd__a2bb2o_2 _34865_ (.A1_N(_01583_),
    .A2_N(_06786_),
    .B1(_04005_),
    .B2(_14593_),
    .X(_06787_));
 sky130_fd_sc_hd__and2_2 _34866_ (.A(_06785_),
    .B(_06787_),
    .X(_06788_));
 sky130_fd_sc_hd__o21ai_2 _34867_ (.A1(_06395_),
    .A2(_06402_),
    .B1(_06788_),
    .Y(_06789_));
 sky130_fd_sc_hd__or3_2 _34868_ (.A(_06395_),
    .B(_06402_),
    .C(_06788_),
    .X(_06790_));
 sky130_fd_sc_hd__nand4_2 _34869_ (.A(_03023_),
    .B(_06783_),
    .C(_06789_),
    .D(_06790_),
    .Y(_06791_));
 sky130_fd_sc_hd__a22o_2 _34870_ (.A1(_03023_),
    .A2(_04905_),
    .B1(_06789_),
    .B2(_06790_),
    .X(_06792_));
 sky130_fd_sc_hd__nand3b_2 _34871_ (.A_N(_06405_),
    .B(_06791_),
    .C(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__a21bo_2 _34872_ (.A1(_06791_),
    .A2(_06792_),
    .B1_N(_06405_),
    .X(_06794_));
 sky130_fd_sc_hd__and2_2 _34873_ (.A(_06430_),
    .B(_06440_),
    .X(_06796_));
 sky130_fd_sc_hd__buf_1 _34874_ (.A(_02643_),
    .X(_06797_));
 sky130_fd_sc_hd__nor2_2 _34875_ (.A(_15155_),
    .B(_06797_),
    .Y(_06798_));
 sky130_fd_sc_hd__o22a_2 _34876_ (.A1(_15155_),
    .A2(_05231_),
    .B1(_06797_),
    .B2(_14949_),
    .X(_06799_));
 sky130_fd_sc_hd__a21o_2 _34877_ (.A1(_06432_),
    .A2(_06798_),
    .B1(_06799_),
    .X(_06800_));
 sky130_fd_sc_hd__nor2_2 _34878_ (.A(_05521_),
    .B(_04187_),
    .Y(_06801_));
 sky130_fd_sc_hd__xnor2_2 _34879_ (.A(_06800_),
    .B(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__xnor2_2 _34880_ (.A(_06393_),
    .B(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__a21oi_2 _34881_ (.A1(_06185_),
    .A2(_06432_),
    .B1(_06435_),
    .Y(_06804_));
 sky130_fd_sc_hd__xnor2_2 _34882_ (.A(_06803_),
    .B(_06804_),
    .Y(_06805_));
 sky130_fd_sc_hd__o21a_2 _34883_ (.A1(_06438_),
    .A2(_06796_),
    .B1(_06805_),
    .X(_06807_));
 sky130_fd_sc_hd__nor3_2 _34884_ (.A(_06438_),
    .B(_06796_),
    .C(_06805_),
    .Y(_06808_));
 sky130_fd_sc_hd__nor2_2 _34885_ (.A(_06807_),
    .B(_06808_),
    .Y(_06809_));
 sky130_fd_sc_hd__or4_2 _34886_ (.A(_05980_),
    .B(_17409_),
    .C(_05504_),
    .D(_05522_),
    .X(_06810_));
 sky130_fd_sc_hd__a22o_2 _34887_ (.A1(_02984_),
    .A2(_00662_),
    .B1(_04138_),
    .B2(_06414_),
    .X(_06811_));
 sky130_fd_sc_hd__and2_2 _34888_ (.A(_06810_),
    .B(_06811_),
    .X(_06812_));
 sky130_fd_sc_hd__buf_1 _34889_ (.A(_03345_),
    .X(_06813_));
 sky130_fd_sc_hd__nand2_2 _34890_ (.A(_06813_),
    .B(_03973_),
    .Y(_06814_));
 sky130_fd_sc_hd__xor2_2 _34891_ (.A(_06812_),
    .B(_06814_),
    .X(_06815_));
 sky130_fd_sc_hd__buf_1 _34892_ (.A(_04162_),
    .X(_06816_));
 sky130_fd_sc_hd__or3b_2 _34893_ (.A(_01804_),
    .B(_01866_),
    .C_N(_06419_),
    .X(_06818_));
 sky130_fd_sc_hd__a21o_2 _34894_ (.A1(_16934_),
    .A2(_03438_),
    .B1(_06419_),
    .X(_06819_));
 sky130_fd_sc_hd__and2_2 _34895_ (.A(_06818_),
    .B(_06819_),
    .X(_06820_));
 sky130_fd_sc_hd__or3b_2 _34896_ (.A(_04847_),
    .B(_06816_),
    .C_N(_06820_),
    .X(_06821_));
 sky130_fd_sc_hd__buf_1 _34897_ (.A(_01862_),
    .X(_06822_));
 sky130_fd_sc_hd__a21o_2 _34898_ (.A1(_16614_),
    .A2(_06822_),
    .B1(_06820_),
    .X(_06823_));
 sky130_fd_sc_hd__nand2_2 _34899_ (.A(_06821_),
    .B(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__nand2_2 _34900_ (.A(_06169_),
    .B(_06419_),
    .Y(_06825_));
 sky130_fd_sc_hd__a21bo_2 _34901_ (.A1(_06421_),
    .A2(_06422_),
    .B1_N(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__xor2_2 _34902_ (.A(_06824_),
    .B(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__nor2_2 _34903_ (.A(_06815_),
    .B(_06827_),
    .Y(_06829_));
 sky130_fd_sc_hd__and2_2 _34904_ (.A(_06815_),
    .B(_06827_),
    .X(_06830_));
 sky130_fd_sc_hd__nor2_2 _34905_ (.A(_06829_),
    .B(_06830_),
    .Y(_06831_));
 sky130_fd_sc_hd__xnor2_2 _34906_ (.A(_06809_),
    .B(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__or2b_2 _34907_ (.A(_06441_),
    .B_N(_06442_),
    .X(_06833_));
 sky130_fd_sc_hd__o21ai_2 _34908_ (.A1(_06429_),
    .A2(_06443_),
    .B1(_06833_),
    .Y(_06834_));
 sky130_fd_sc_hd__xnor2_2 _34909_ (.A(_06832_),
    .B(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__nand3_2 _34910_ (.A(_06793_),
    .B(_06794_),
    .C(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__a21o_2 _34911_ (.A1(_06793_),
    .A2(_06794_),
    .B1(_06835_),
    .X(_06837_));
 sky130_fd_sc_hd__o211a_2 _34912_ (.A1(_06407_),
    .A2(_06450_),
    .B1(_06836_),
    .C1(_06837_),
    .X(_06838_));
 sky130_fd_sc_hd__a211oi_2 _34913_ (.A1(_06836_),
    .A2(_06837_),
    .B1(_06407_),
    .C1(_06450_),
    .Y(_06840_));
 sky130_fd_sc_hd__o21ai_2 _34914_ (.A1(_06501_),
    .A2(_06502_),
    .B1(_06499_),
    .Y(_06841_));
 sky130_fd_sc_hd__or2b_2 _34915_ (.A(_06480_),
    .B_N(_06504_),
    .X(_06842_));
 sky130_fd_sc_hd__nand2_2 _34916_ (.A(_06841_),
    .B(_06842_),
    .Y(_06843_));
 sky130_fd_sc_hd__a21o_2 _34917_ (.A1(_06409_),
    .A2(_06448_),
    .B1(_06446_),
    .X(_06844_));
 sky130_fd_sc_hd__o31ai_2 _34918_ (.A1(_01583_),
    .A2(_05441_),
    .A3(_06463_),
    .B1(_06461_),
    .Y(_06845_));
 sky130_fd_sc_hd__or3_2 _34919_ (.A(_03378_),
    .B(_05931_),
    .C(_06460_),
    .X(_06846_));
 sky130_fd_sc_hd__nor2_2 _34920_ (.A(_02471_),
    .B(_05931_),
    .Y(_06847_));
 sky130_fd_sc_hd__a21o_2 _34921_ (.A1(_02989_),
    .A2(_02928_),
    .B1(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__and4_2 _34922_ (.A(_02983_),
    .B(_04451_),
    .C(_06846_),
    .D(_06848_),
    .X(_06849_));
 sky130_fd_sc_hd__o2bb2a_2 _34923_ (.A1_N(_06846_),
    .A2_N(_06848_),
    .B1(_02463_),
    .B2(_03318_),
    .X(_06851_));
 sky130_fd_sc_hd__nor2_2 _34924_ (.A(_06849_),
    .B(_06851_),
    .Y(_06852_));
 sky130_fd_sc_hd__nand2_2 _34925_ (.A(_04837_),
    .B(_00567_),
    .Y(_06853_));
 sky130_fd_sc_hd__a22o_2 _34926_ (.A1(_04837_),
    .A2(_05450_),
    .B1(_00567_),
    .B2(_01040_),
    .X(_06854_));
 sky130_fd_sc_hd__o21ai_2 _34927_ (.A1(_06466_),
    .A2(_06853_),
    .B1(_06854_),
    .Y(_06855_));
 sky130_fd_sc_hd__nand2_2 _34928_ (.A(_00633_),
    .B(_03327_),
    .Y(_06856_));
 sky130_fd_sc_hd__xnor2_2 _34929_ (.A(_06855_),
    .B(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__or2_2 _34930_ (.A(_06468_),
    .B(_06469_),
    .X(_06858_));
 sky130_fd_sc_hd__o21a_2 _34931_ (.A1(_06102_),
    .A2(_06466_),
    .B1(_06858_),
    .X(_06859_));
 sky130_fd_sc_hd__nor2_2 _34932_ (.A(_06857_),
    .B(_06859_),
    .Y(_06860_));
 sky130_fd_sc_hd__and2_2 _34933_ (.A(_06857_),
    .B(_06859_),
    .X(_06862_));
 sky130_fd_sc_hd__nor2_2 _34934_ (.A(_06860_),
    .B(_06862_),
    .Y(_06863_));
 sky130_fd_sc_hd__xnor2_2 _34935_ (.A(_06852_),
    .B(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__a21o_2 _34936_ (.A1(_06465_),
    .A2(_06473_),
    .B1(_06472_),
    .X(_06865_));
 sky130_fd_sc_hd__xnor2_2 _34937_ (.A(_06864_),
    .B(_06865_),
    .Y(_06866_));
 sky130_fd_sc_hd__xnor2_2 _34938_ (.A(_06845_),
    .B(_06866_),
    .Y(_06867_));
 sky130_fd_sc_hd__or2b_2 _34939_ (.A(_06495_),
    .B_N(_06487_),
    .X(_06868_));
 sky130_fd_sc_hd__a21bo_2 _34940_ (.A1(_06485_),
    .A2(_06496_),
    .B1_N(_06868_),
    .X(_06869_));
 sky130_fd_sc_hd__o21a_2 _34941_ (.A1(_06418_),
    .A2(_06428_),
    .B1(_06426_),
    .X(_06870_));
 sky130_fd_sc_hd__a31o_2 _34942_ (.A1(_04837_),
    .A2(_06484_),
    .A3(_06493_),
    .B1(_06490_),
    .X(_06871_));
 sky130_fd_sc_hd__a21bo_2 _34943_ (.A1(_06415_),
    .A2(_06417_),
    .B1_N(_06410_),
    .X(_06873_));
 sky130_fd_sc_hd__and4_2 _34944_ (.A(_03024_),
    .B(_05507_),
    .C(_18328_),
    .D(_06488_),
    .X(_06874_));
 sky130_fd_sc_hd__o22a_2 _34945_ (.A1(_05979_),
    .A2(_06491_),
    .B1(_18344_),
    .B2(_04501_),
    .X(_06875_));
 sky130_fd_sc_hd__nor2_2 _34946_ (.A(_06874_),
    .B(_06875_),
    .Y(_06876_));
 sky130_fd_sc_hd__nand2_2 _34947_ (.A(_01837_),
    .B(_04469_),
    .Y(_06877_));
 sky130_fd_sc_hd__xor2_2 _34948_ (.A(_06876_),
    .B(_06877_),
    .X(_06878_));
 sky130_fd_sc_hd__xnor2_2 _34949_ (.A(_06873_),
    .B(_06878_),
    .Y(_06879_));
 sky130_fd_sc_hd__xnor2_2 _34950_ (.A(_06871_),
    .B(_06879_),
    .Y(_06880_));
 sky130_fd_sc_hd__xnor2_2 _34951_ (.A(_06870_),
    .B(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__xnor2_2 _34952_ (.A(_06869_),
    .B(_06881_),
    .Y(_06882_));
 sky130_fd_sc_hd__nor2_2 _34953_ (.A(_06483_),
    .B(_06497_),
    .Y(_06884_));
 sky130_fd_sc_hd__and2b_2 _34954_ (.A_N(_06498_),
    .B(_06482_),
    .X(_06885_));
 sky130_fd_sc_hd__nor2_2 _34955_ (.A(_06884_),
    .B(_06885_),
    .Y(_06886_));
 sky130_fd_sc_hd__xnor2_2 _34956_ (.A(_06882_),
    .B(_06886_),
    .Y(_06887_));
 sky130_fd_sc_hd__xnor2_2 _34957_ (.A(_06867_),
    .B(_06887_),
    .Y(_06888_));
 sky130_fd_sc_hd__xnor2_2 _34958_ (.A(_06844_),
    .B(_06888_),
    .Y(_06889_));
 sky130_fd_sc_hd__xor2_2 _34959_ (.A(_06843_),
    .B(_06889_),
    .X(_06890_));
 sky130_fd_sc_hd__or3_2 _34960_ (.A(_06838_),
    .B(_06840_),
    .C(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__o21ai_2 _34961_ (.A1(_06838_),
    .A2(_06840_),
    .B1(_06890_),
    .Y(_06892_));
 sky130_fd_sc_hd__o211a_2 _34962_ (.A1(_06452_),
    .A2(_06782_),
    .B1(_06891_),
    .C1(_06892_),
    .X(_06893_));
 sky130_fd_sc_hd__a211oi_2 _34963_ (.A1(_06891_),
    .A2(_06892_),
    .B1(_06452_),
    .C1(_06782_),
    .Y(_06895_));
 sky130_fd_sc_hd__and2b_2 _34964_ (.A_N(_06506_),
    .B(_06457_),
    .X(_06896_));
 sky130_fd_sc_hd__a21oi_2 _34965_ (.A1(_06458_),
    .A2(_06505_),
    .B1(_06896_),
    .Y(_06897_));
 sky130_fd_sc_hd__a21oi_2 _34966_ (.A1(_06459_),
    .A2(_06479_),
    .B1(_06476_),
    .Y(_06898_));
 sky130_fd_sc_hd__xnor2_2 _34967_ (.A(_06897_),
    .B(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__or3_2 _34968_ (.A(_06893_),
    .B(_06895_),
    .C(_06899_),
    .X(_06900_));
 sky130_fd_sc_hd__o21ai_2 _34969_ (.A1(_06893_),
    .A2(_06895_),
    .B1(_06899_),
    .Y(_06901_));
 sky130_fd_sc_hd__o211ai_2 _34970_ (.A1(_06510_),
    .A2(_06519_),
    .B1(_06900_),
    .C1(_06901_),
    .Y(_06902_));
 sky130_fd_sc_hd__a211o_2 _34971_ (.A1(_06900_),
    .A2(_06901_),
    .B1(_06510_),
    .C1(_06519_),
    .X(_06903_));
 sky130_fd_sc_hd__and3_2 _34972_ (.A(_06516_),
    .B(_06902_),
    .C(_06903_),
    .X(_06904_));
 sky130_fd_sc_hd__a21oi_2 _34973_ (.A1(_06902_),
    .A2(_06903_),
    .B1(_06516_),
    .Y(_06906_));
 sky130_fd_sc_hd__a211o_2 _34974_ (.A1(_06521_),
    .A2(_06781_),
    .B1(_06904_),
    .C1(_06906_),
    .X(_06907_));
 sky130_fd_sc_hd__o211ai_2 _34975_ (.A1(_06904_),
    .A2(_06906_),
    .B1(_06521_),
    .C1(_06781_),
    .Y(_06908_));
 sky130_fd_sc_hd__nand2_2 _34976_ (.A(_06907_),
    .B(_06908_),
    .Y(_06909_));
 sky130_fd_sc_hd__inv_2 _34977_ (.A(_06060_),
    .Y(_06910_));
 sky130_fd_sc_hd__or3_2 _34978_ (.A(_06221_),
    .B(_06526_),
    .C(_06527_),
    .X(_06911_));
 sky130_fd_sc_hd__a2111o_2 _34979_ (.A1(_05421_),
    .A2(_05425_),
    .B1(_06910_),
    .C1(_06911_),
    .D1(_05588_),
    .X(_06912_));
 sky130_fd_sc_hd__or2_2 _34980_ (.A(_06380_),
    .B(_06527_),
    .X(_06913_));
 sky130_fd_sc_hd__bufinv_8 _34981_ (.A(_06526_),
    .Y(_06914_));
 sky130_fd_sc_hd__o211a_2 _34982_ (.A1(_06224_),
    .A2(_06911_),
    .B1(_06913_),
    .C1(_06914_),
    .X(_06915_));
 sky130_fd_sc_hd__nand2_2 _34983_ (.A(_06912_),
    .B(_06915_),
    .Y(_06917_));
 sky130_fd_sc_hd__xnor2_2 _34984_ (.A(_06909_),
    .B(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__and2b_2 _34985_ (.A_N(_06780_),
    .B(_06918_),
    .X(_06919_));
 sky130_fd_sc_hd__nor2b_2 _34986_ (.A(_06918_),
    .B_N(_06780_),
    .Y(_06920_));
 sky130_fd_sc_hd__nor2_2 _34987_ (.A(_06919_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__xnor2_2 _34988_ (.A(_14335_),
    .B(_06921_),
    .Y(_06922_));
 sky130_fd_sc_hd__and2b_2 _34989_ (.A_N(_06529_),
    .B(_06650_),
    .X(_06923_));
 sky130_fd_sc_hd__a21oi_2 _34990_ (.A1(_14204_),
    .A2(_06651_),
    .B1(_06923_),
    .Y(_06924_));
 sky130_fd_sc_hd__xnor2_2 _34991_ (.A(_06922_),
    .B(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__inv_2 _34992_ (.A(_06653_),
    .Y(_06926_));
 sky130_fd_sc_hd__o21a_2 _34993_ (.A1(_06378_),
    .A2(_06652_),
    .B1(_06361_),
    .X(_06928_));
 sky130_fd_sc_hd__a21oi_2 _34994_ (.A1(_06378_),
    .A2(_06652_),
    .B1(_06928_),
    .Y(_06929_));
 sky130_fd_sc_hd__o31a_2 _34995_ (.A1(_06375_),
    .A2(_06370_),
    .A3(_06926_),
    .B1(_06929_),
    .X(_06930_));
 sky130_fd_sc_hd__or2_2 _34996_ (.A(_06925_),
    .B(_06930_),
    .X(_06931_));
 sky130_fd_sc_hd__nand2_2 _34997_ (.A(_06925_),
    .B(_06930_),
    .Y(_06932_));
 sky130_fd_sc_hd__nand2_2 _34998_ (.A(_06931_),
    .B(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__nor2_2 _34999_ (.A(_14499_),
    .B(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__and2_2 _35000_ (.A(_14499_),
    .B(_06933_),
    .X(_06935_));
 sky130_fd_sc_hd__nor2_2 _35001_ (.A(_06934_),
    .B(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__o21ba_2 _35002_ (.A1(_06659_),
    .A2(_06657_),
    .B1_N(_06656_),
    .X(_06937_));
 sky130_fd_sc_hd__a21oi_2 _35003_ (.A1(_06373_),
    .A2(_06658_),
    .B1(_06937_),
    .Y(_06939_));
 sky130_fd_sc_hd__xnor2_2 _35004_ (.A(_06936_),
    .B(_06939_),
    .Y(oO[76]));
 sky130_fd_sc_hd__or2_2 _35005_ (.A(_06922_),
    .B(_06924_),
    .X(_06940_));
 sky130_fd_sc_hd__a21o_2 _35006_ (.A1(_06912_),
    .A2(_06915_),
    .B1(_06909_),
    .X(_06941_));
 sky130_fd_sc_hd__nor2_2 _35007_ (.A(_06897_),
    .B(_06898_),
    .Y(_06942_));
 sky130_fd_sc_hd__nor3_2 _35008_ (.A(_06893_),
    .B(_06895_),
    .C(_06899_),
    .Y(_06943_));
 sky130_fd_sc_hd__inv_2 _35009_ (.A(_06838_),
    .Y(_06944_));
 sky130_fd_sc_hd__and3b_2 _35010_ (.A_N(_06405_),
    .B(_06791_),
    .C(_06792_),
    .X(_06945_));
 sky130_fd_sc_hd__and3_2 _35011_ (.A(_06793_),
    .B(_06794_),
    .C(_06835_),
    .X(_06946_));
 sky130_fd_sc_hd__o22a_2 _35012_ (.A1(_02463_),
    .A2(_06786_),
    .B1(_04901_),
    .B2(_01028_),
    .X(_06947_));
 sky130_fd_sc_hd__or2_2 _35013_ (.A(_00228_),
    .B(_06399_),
    .X(_06949_));
 sky130_fd_sc_hd__and2b_2 _35014_ (.A_N(_06947_),
    .B(_06949_),
    .X(_06950_));
 sky130_fd_sc_hd__nand3_2 _35015_ (.A(_06785_),
    .B(_06789_),
    .C(_06950_),
    .Y(_06951_));
 sky130_fd_sc_hd__a21o_2 _35016_ (.A1(_06785_),
    .A2(_06789_),
    .B1(_06950_),
    .X(_06952_));
 sky130_fd_sc_hd__a21o_2 _35017_ (.A1(_06951_),
    .A2(_06952_),
    .B1(_06791_),
    .X(_06953_));
 sky130_fd_sc_hd__nand3_2 _35018_ (.A(_06791_),
    .B(_06951_),
    .C(_06952_),
    .Y(_06954_));
 sky130_fd_sc_hd__and3_2 _35019_ (.A(_01033_),
    .B(_03454_),
    .C(_06798_),
    .X(_06955_));
 sky130_fd_sc_hd__a21oi_2 _35020_ (.A1(_01033_),
    .A2(_03454_),
    .B1(_06798_),
    .Y(_06956_));
 sky130_fd_sc_hd__nor2_2 _35021_ (.A(_06955_),
    .B(_06956_),
    .Y(_06957_));
 sky130_fd_sc_hd__nor2_2 _35022_ (.A(_05521_),
    .B(_05231_),
    .Y(_06958_));
 sky130_fd_sc_hd__xnor2_2 _35023_ (.A(_06957_),
    .B(_06958_),
    .Y(_06960_));
 sky130_fd_sc_hd__nand2_2 _35024_ (.A(_06432_),
    .B(_06798_),
    .Y(_06961_));
 sky130_fd_sc_hd__o31a_2 _35025_ (.A1(_05521_),
    .A2(_04187_),
    .A3(_06799_),
    .B1(_06961_),
    .X(_06962_));
 sky130_fd_sc_hd__nor2_2 _35026_ (.A(_06960_),
    .B(_06962_),
    .Y(_06963_));
 sky130_fd_sc_hd__and2_2 _35027_ (.A(_06960_),
    .B(_06962_),
    .X(_06964_));
 sky130_fd_sc_hd__or2_2 _35028_ (.A(_06963_),
    .B(_06964_),
    .X(_06965_));
 sky130_fd_sc_hd__inv_2 _35029_ (.A(_06802_),
    .Y(_06966_));
 sky130_fd_sc_hd__or2b_2 _35030_ (.A(_06804_),
    .B_N(_06803_),
    .X(_06967_));
 sky130_fd_sc_hd__o21a_2 _35031_ (.A1(_06393_),
    .A2(_06966_),
    .B1(_06967_),
    .X(_06968_));
 sky130_fd_sc_hd__or2_2 _35032_ (.A(_06965_),
    .B(_06968_),
    .X(_06969_));
 sky130_fd_sc_hd__nand2_2 _35033_ (.A(_06965_),
    .B(_06968_),
    .Y(_06971_));
 sky130_fd_sc_hd__and2_2 _35034_ (.A(_06969_),
    .B(_06971_),
    .X(_06972_));
 sky130_fd_sc_hd__or4_2 _35035_ (.A(_05980_),
    .B(_05978_),
    .C(_05522_),
    .D(_06816_),
    .X(_06973_));
 sky130_fd_sc_hd__a22o_2 _35036_ (.A1(_06411_),
    .A2(_04138_),
    .B1(_06822_),
    .B2(_06414_),
    .X(_06974_));
 sky130_fd_sc_hd__a22o_2 _35037_ (.A1(_06813_),
    .A2(_06413_),
    .B1(_06973_),
    .B2(_06974_),
    .X(_06975_));
 sky130_fd_sc_hd__nand4_2 _35038_ (.A(_06813_),
    .B(_06413_),
    .C(_06973_),
    .D(_06974_),
    .Y(_06976_));
 sky130_fd_sc_hd__nand2_2 _35039_ (.A(_06975_),
    .B(_06976_),
    .Y(_06977_));
 sky130_fd_sc_hd__or2_2 _35040_ (.A(_16606_),
    .B(_04187_),
    .X(_06978_));
 sky130_fd_sc_hd__or3_2 _35041_ (.A(_01804_),
    .B(_05543_),
    .C(_06978_),
    .X(_06979_));
 sky130_fd_sc_hd__a2bb2o_2 _35042_ (.A1_N(_16606_),
    .A2_N(_05543_),
    .B1(_02648_),
    .B2(_16934_),
    .X(_06980_));
 sky130_fd_sc_hd__nand2_2 _35043_ (.A(_06979_),
    .B(_06980_),
    .Y(_06982_));
 sky130_fd_sc_hd__buf_1 _35044_ (.A(_02629_),
    .X(_06983_));
 sky130_fd_sc_hd__nand2_2 _35045_ (.A(_16614_),
    .B(_06983_),
    .Y(_06984_));
 sky130_fd_sc_hd__xnor2_2 _35046_ (.A(_06982_),
    .B(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__a21o_2 _35047_ (.A1(_06818_),
    .A2(_06821_),
    .B1(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__nand3_2 _35048_ (.A(_06818_),
    .B(_06821_),
    .C(_06985_),
    .Y(_06987_));
 sky130_fd_sc_hd__nand2_2 _35049_ (.A(_06986_),
    .B(_06987_),
    .Y(_06988_));
 sky130_fd_sc_hd__xor2_2 _35050_ (.A(_06977_),
    .B(_06988_),
    .X(_06989_));
 sky130_fd_sc_hd__nand2_2 _35051_ (.A(_06972_),
    .B(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__or2_2 _35052_ (.A(_06972_),
    .B(_06989_),
    .X(_06991_));
 sky130_fd_sc_hd__nand2_2 _35053_ (.A(_06990_),
    .B(_06991_),
    .Y(_06993_));
 sky130_fd_sc_hd__a21oi_2 _35054_ (.A1(_06809_),
    .A2(_06831_),
    .B1(_06807_),
    .Y(_06994_));
 sky130_fd_sc_hd__nor2_2 _35055_ (.A(_06993_),
    .B(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__and2_2 _35056_ (.A(_06993_),
    .B(_06994_),
    .X(_06996_));
 sky130_fd_sc_hd__nor2_2 _35057_ (.A(_06995_),
    .B(_06996_),
    .Y(_06997_));
 sky130_fd_sc_hd__nand3_2 _35058_ (.A(_06953_),
    .B(_06954_),
    .C(_06997_),
    .Y(_06998_));
 sky130_fd_sc_hd__a21o_2 _35059_ (.A1(_06953_),
    .A2(_06954_),
    .B1(_06997_),
    .X(_06999_));
 sky130_fd_sc_hd__o211ai_2 _35060_ (.A1(_06945_),
    .A2(_06946_),
    .B1(_06998_),
    .C1(_06999_),
    .Y(_07000_));
 sky130_fd_sc_hd__a211o_2 _35061_ (.A1(_06998_),
    .A2(_06999_),
    .B1(_06945_),
    .C1(_06946_),
    .X(_07001_));
 sky130_fd_sc_hd__o21ai_2 _35062_ (.A1(_06884_),
    .A2(_06885_),
    .B1(_06882_),
    .Y(_07002_));
 sky130_fd_sc_hd__or2b_2 _35063_ (.A(_06867_),
    .B_N(_06887_),
    .X(_07004_));
 sky130_fd_sc_hd__nand2_2 _35064_ (.A(_07002_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__and2b_2 _35065_ (.A_N(_06832_),
    .B(_06834_),
    .X(_07006_));
 sky130_fd_sc_hd__buf_1 _35066_ (.A(_04781_),
    .X(_07007_));
 sky130_fd_sc_hd__a31o_2 _35067_ (.A1(_02989_),
    .A2(_07007_),
    .A3(_06847_),
    .B1(_06849_),
    .X(_07008_));
 sky130_fd_sc_hd__nand2_2 _35068_ (.A(_00633_),
    .B(_02928_),
    .Y(_07009_));
 sky130_fd_sc_hd__or3_2 _35069_ (.A(_03378_),
    .B(_05931_),
    .C(_07009_),
    .X(_07010_));
 sky130_fd_sc_hd__o21ai_2 _35070_ (.A1(_03378_),
    .A2(_05931_),
    .B1(_07009_),
    .Y(_07011_));
 sky130_fd_sc_hd__nand2_2 _35071_ (.A(_07010_),
    .B(_07011_),
    .Y(_07012_));
 sky130_fd_sc_hd__nor2_2 _35072_ (.A(_02471_),
    .B(_03318_),
    .Y(_07013_));
 sky130_fd_sc_hd__xnor2_2 _35073_ (.A(_07012_),
    .B(_07013_),
    .Y(_07015_));
 sky130_fd_sc_hd__nand2_2 _35074_ (.A(_01837_),
    .B(_05450_),
    .Y(_07016_));
 sky130_fd_sc_hd__xnor2_2 _35075_ (.A(_06853_),
    .B(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__or3_2 _35076_ (.A(_03389_),
    .B(_00944_),
    .C(_07017_),
    .X(_07018_));
 sky130_fd_sc_hd__o21ai_2 _35077_ (.A1(_03389_),
    .A2(_00944_),
    .B1(_07017_),
    .Y(_07019_));
 sky130_fd_sc_hd__nand2_2 _35078_ (.A(_07018_),
    .B(_07019_),
    .Y(_07020_));
 sky130_fd_sc_hd__o22a_2 _35079_ (.A1(_06466_),
    .A2(_06853_),
    .B1(_06855_),
    .B2(_06856_),
    .X(_07021_));
 sky130_fd_sc_hd__nor2_2 _35080_ (.A(_07020_),
    .B(_07021_),
    .Y(_07022_));
 sky130_fd_sc_hd__nand2_2 _35081_ (.A(_07020_),
    .B(_07021_),
    .Y(_07023_));
 sky130_fd_sc_hd__and2b_2 _35082_ (.A_N(_07022_),
    .B(_07023_),
    .X(_07024_));
 sky130_fd_sc_hd__xnor2_2 _35083_ (.A(_07015_),
    .B(_07024_),
    .Y(_07026_));
 sky130_fd_sc_hd__a21o_2 _35084_ (.A1(_06852_),
    .A2(_06863_),
    .B1(_06860_),
    .X(_07027_));
 sky130_fd_sc_hd__xnor2_2 _35085_ (.A(_07026_),
    .B(_07027_),
    .Y(_07028_));
 sky130_fd_sc_hd__xnor2_2 _35086_ (.A(_07008_),
    .B(_07028_),
    .Y(_07029_));
 sky130_fd_sc_hd__nor2_2 _35087_ (.A(_06870_),
    .B(_06880_),
    .Y(_07030_));
 sky130_fd_sc_hd__and2b_2 _35088_ (.A_N(_06881_),
    .B(_06869_),
    .X(_07031_));
 sky130_fd_sc_hd__or2b_2 _35089_ (.A(_06878_),
    .B_N(_06873_),
    .X(_07032_));
 sky130_fd_sc_hd__a21bo_2 _35090_ (.A1(_06871_),
    .A2(_06879_),
    .B1_N(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__a31o_2 _35091_ (.A1(_06821_),
    .A2(_06823_),
    .A3(_06826_),
    .B1(_06829_),
    .X(_07034_));
 sky130_fd_sc_hd__a31o_2 _35092_ (.A1(_01837_),
    .A2(_06484_),
    .A3(_06876_),
    .B1(_06874_),
    .X(_07035_));
 sky130_fd_sc_hd__or3b_2 _35093_ (.A(_05500_),
    .B(_04862_),
    .C_N(_06812_),
    .X(_07037_));
 sky130_fd_sc_hd__nand2_2 _35094_ (.A(_06810_),
    .B(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__buf_1 _35095_ (.A(_18328_),
    .X(_07039_));
 sky130_fd_sc_hd__and4_2 _35096_ (.A(_05507_),
    .B(_03973_),
    .C(_07039_),
    .D(_06488_),
    .X(_07040_));
 sky130_fd_sc_hd__o22a_2 _35097_ (.A1(_04862_),
    .A2(_06491_),
    .B1(_18344_),
    .B2(_05979_),
    .X(_07041_));
 sky130_fd_sc_hd__nor2_2 _35098_ (.A(_07040_),
    .B(_07041_),
    .Y(_07042_));
 sky130_fd_sc_hd__nand2_2 _35099_ (.A(_03024_),
    .B(_04469_),
    .Y(_07043_));
 sky130_fd_sc_hd__xor2_2 _35100_ (.A(_07042_),
    .B(_07043_),
    .X(_07044_));
 sky130_fd_sc_hd__xnor2_2 _35101_ (.A(_07038_),
    .B(_07044_),
    .Y(_07045_));
 sky130_fd_sc_hd__xnor2_2 _35102_ (.A(_07035_),
    .B(_07045_),
    .Y(_07046_));
 sky130_fd_sc_hd__xnor2_2 _35103_ (.A(_07034_),
    .B(_07046_),
    .Y(_07048_));
 sky130_fd_sc_hd__xor2_2 _35104_ (.A(_07033_),
    .B(_07048_),
    .X(_07049_));
 sky130_fd_sc_hd__o21a_2 _35105_ (.A1(_07030_),
    .A2(_07031_),
    .B1(_07049_),
    .X(_07050_));
 sky130_fd_sc_hd__nor3_2 _35106_ (.A(_07030_),
    .B(_07031_),
    .C(_07049_),
    .Y(_07051_));
 sky130_fd_sc_hd__nor2_2 _35107_ (.A(_07050_),
    .B(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__xnor2_2 _35108_ (.A(_07029_),
    .B(_07052_),
    .Y(_07053_));
 sky130_fd_sc_hd__xnor2_2 _35109_ (.A(_07006_),
    .B(_07053_),
    .Y(_07054_));
 sky130_fd_sc_hd__xnor2_2 _35110_ (.A(_07005_),
    .B(_07054_),
    .Y(_07055_));
 sky130_fd_sc_hd__and3_2 _35111_ (.A(_07000_),
    .B(_07001_),
    .C(_07055_),
    .X(_07056_));
 sky130_fd_sc_hd__a21oi_2 _35112_ (.A1(_07000_),
    .A2(_07001_),
    .B1(_07055_),
    .Y(_07057_));
 sky130_fd_sc_hd__a211o_2 _35113_ (.A1(_06944_),
    .A2(_06891_),
    .B1(_07056_),
    .C1(_07057_),
    .X(_07059_));
 sky130_fd_sc_hd__o211ai_2 _35114_ (.A1(_07056_),
    .A2(_07057_),
    .B1(_06944_),
    .C1(_06891_),
    .Y(_07060_));
 sky130_fd_sc_hd__nand2_2 _35115_ (.A(_06844_),
    .B(_06888_),
    .Y(_07061_));
 sky130_fd_sc_hd__or2b_2 _35116_ (.A(_06889_),
    .B_N(_06843_),
    .X(_07062_));
 sky130_fd_sc_hd__and2b_2 _35117_ (.A_N(_06864_),
    .B(_06865_),
    .X(_07063_));
 sky130_fd_sc_hd__a21oi_2 _35118_ (.A1(_06845_),
    .A2(_06866_),
    .B1(_07063_),
    .Y(_07064_));
 sky130_fd_sc_hd__a21o_2 _35119_ (.A1(_07061_),
    .A2(_07062_),
    .B1(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__nand3_2 _35120_ (.A(_07061_),
    .B(_07062_),
    .C(_07064_),
    .Y(_07066_));
 sky130_fd_sc_hd__and2_2 _35121_ (.A(_07065_),
    .B(_07066_),
    .X(_07067_));
 sky130_fd_sc_hd__nand3_2 _35122_ (.A(_07059_),
    .B(_07060_),
    .C(_07067_),
    .Y(_07068_));
 sky130_fd_sc_hd__a21o_2 _35123_ (.A1(_07059_),
    .A2(_07060_),
    .B1(_07067_),
    .X(_07070_));
 sky130_fd_sc_hd__o211ai_2 _35124_ (.A1(_06893_),
    .A2(_06943_),
    .B1(_07068_),
    .C1(_07070_),
    .Y(_07071_));
 sky130_fd_sc_hd__a211o_2 _35125_ (.A1(_07068_),
    .A2(_07070_),
    .B1(_06893_),
    .C1(_06943_),
    .X(_07072_));
 sky130_fd_sc_hd__and3_2 _35126_ (.A(_06942_),
    .B(_07071_),
    .C(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__a21oi_2 _35127_ (.A1(_07071_),
    .A2(_07072_),
    .B1(_06942_),
    .Y(_07074_));
 sky130_fd_sc_hd__or2_2 _35128_ (.A(_07073_),
    .B(_07074_),
    .X(_07075_));
 sky130_fd_sc_hd__a21boi_2 _35129_ (.A1(_06516_),
    .A2(_06903_),
    .B1_N(_06902_),
    .Y(_07076_));
 sky130_fd_sc_hd__xor2_2 _35130_ (.A(_07075_),
    .B(_07076_),
    .X(_07077_));
 sky130_fd_sc_hd__nand3_2 _35131_ (.A(_06907_),
    .B(_06941_),
    .C(_07077_),
    .Y(_07078_));
 sky130_fd_sc_hd__a21o_2 _35132_ (.A1(_06907_),
    .A2(_06941_),
    .B1(_07077_),
    .X(_07079_));
 sky130_fd_sc_hd__and2b_2 _35133_ (.A_N(_06760_),
    .B(_06761_),
    .X(_07081_));
 sky130_fd_sc_hd__nand2_2 _35134_ (.A(_06707_),
    .B(_06750_),
    .Y(_07082_));
 sky130_fd_sc_hd__nand2_2 _35135_ (.A(iY[46]),
    .B(iX[63]),
    .Y(_07083_));
 sky130_fd_sc_hd__a21o_2 _35136_ (.A1(_06567_),
    .A2(_06681_),
    .B1(_06692_),
    .X(_07084_));
 sky130_fd_sc_hd__nand2_2 _35137_ (.A(_06682_),
    .B(_06691_),
    .Y(_07085_));
 sky130_fd_sc_hd__and2_2 _35138_ (.A(iY[48]),
    .B(iX[62]),
    .X(_07086_));
 sky130_fd_sc_hd__and3_2 _35139_ (.A(iY[47]),
    .B(iX[61]),
    .C(_07086_),
    .X(_07087_));
 sky130_fd_sc_hd__a22oi_2 _35140_ (.A1(iY[48]),
    .A2(iX[61]),
    .B1(iX[62]),
    .B2(iY[47]),
    .Y(_07088_));
 sky130_fd_sc_hd__nor2_2 _35141_ (.A(_07087_),
    .B(_07088_),
    .Y(_07089_));
 sky130_fd_sc_hd__nand2_2 _35142_ (.A(iY[49]),
    .B(iX[60]),
    .Y(_07090_));
 sky130_fd_sc_hd__xnor2_2 _35143_ (.A(_07089_),
    .B(_07090_),
    .Y(_07092_));
 sky130_fd_sc_hd__and2_2 _35144_ (.A(_06662_),
    .B(_07092_),
    .X(_07093_));
 sky130_fd_sc_hd__nor2_2 _35145_ (.A(_06662_),
    .B(_07092_),
    .Y(_07094_));
 sky130_fd_sc_hd__or2_2 _35146_ (.A(_07093_),
    .B(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__a31o_2 _35147_ (.A1(iY[49]),
    .A2(iX[59]),
    .A3(_06685_),
    .B1(_06683_),
    .X(_07096_));
 sky130_fd_sc_hd__and2b_2 _35148_ (.A_N(_07095_),
    .B(_07096_),
    .X(_07097_));
 sky130_fd_sc_hd__and2b_2 _35149_ (.A_N(_07096_),
    .B(_07095_),
    .X(_07098_));
 sky130_fd_sc_hd__or2_2 _35150_ (.A(_07097_),
    .B(_07098_),
    .X(_07099_));
 sky130_fd_sc_hd__a21oi_2 _35151_ (.A1(_06689_),
    .A2(_07085_),
    .B1(_07099_),
    .Y(_07100_));
 sky130_fd_sc_hd__and3_2 _35152_ (.A(_06689_),
    .B(_07085_),
    .C(_07099_),
    .X(_07101_));
 sky130_fd_sc_hd__and4_2 _35153_ (.A(iY[53]),
    .B(iY[54]),
    .C(iX[55]),
    .D(iX[56]),
    .X(_07103_));
 sky130_fd_sc_hd__a22oi_2 _35154_ (.A1(iY[54]),
    .A2(iX[55]),
    .B1(iX[56]),
    .B2(iY[53]),
    .Y(_07104_));
 sky130_fd_sc_hd__nor2_2 _35155_ (.A(_07103_),
    .B(_07104_),
    .Y(_07105_));
 sky130_fd_sc_hd__nand2_2 _35156_ (.A(iX[54]),
    .B(iY[55]),
    .Y(_07106_));
 sky130_fd_sc_hd__xnor2_2 _35157_ (.A(_07105_),
    .B(_07106_),
    .Y(_07107_));
 sky130_fd_sc_hd__and4_2 _35158_ (.A(iY[50]),
    .B(iY[51]),
    .C(iX[58]),
    .D(iX[59]),
    .X(_07108_));
 sky130_fd_sc_hd__a22oi_2 _35159_ (.A1(iY[51]),
    .A2(iX[58]),
    .B1(iX[59]),
    .B2(iY[50]),
    .Y(_07109_));
 sky130_fd_sc_hd__nor2_2 _35160_ (.A(_07108_),
    .B(_07109_),
    .Y(_07110_));
 sky130_fd_sc_hd__nand2_2 _35161_ (.A(iY[52]),
    .B(iX[57]),
    .Y(_07111_));
 sky130_fd_sc_hd__xnor2_2 _35162_ (.A(_07110_),
    .B(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__o21ba_2 _35163_ (.A1(_06671_),
    .A2(_06673_),
    .B1_N(_06670_),
    .X(_07114_));
 sky130_fd_sc_hd__xnor2_2 _35164_ (.A(_07112_),
    .B(_07114_),
    .Y(_07115_));
 sky130_fd_sc_hd__and2_2 _35165_ (.A(_07107_),
    .B(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__nor2_2 _35166_ (.A(_07107_),
    .B(_07115_),
    .Y(_07117_));
 sky130_fd_sc_hd__or2_2 _35167_ (.A(_07116_),
    .B(_07117_),
    .X(_07118_));
 sky130_fd_sc_hd__nor3_2 _35168_ (.A(_07100_),
    .B(_07101_),
    .C(_07118_),
    .Y(_07119_));
 sky130_fd_sc_hd__o21a_2 _35169_ (.A1(_07100_),
    .A2(_07101_),
    .B1(_07118_),
    .X(_07120_));
 sky130_fd_sc_hd__a211oi_2 _35170_ (.A1(_07084_),
    .A2(_06695_),
    .B1(_07119_),
    .C1(_07120_),
    .Y(_07121_));
 sky130_fd_sc_hd__o211a_2 _35171_ (.A1(_07119_),
    .A2(_07120_),
    .B1(_07084_),
    .C1(_06695_),
    .X(_07122_));
 sky130_fd_sc_hd__nor2_2 _35172_ (.A(_07121_),
    .B(_07122_),
    .Y(_07123_));
 sky130_fd_sc_hd__xnor2_2 _35173_ (.A(_07083_),
    .B(_07123_),
    .Y(_07125_));
 sky130_fd_sc_hd__xnor2_2 _35174_ (.A(_06702_),
    .B(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__inv_2 _35175_ (.A(_06746_),
    .Y(_07127_));
 sky130_fd_sc_hd__or2b_2 _35176_ (.A(_06714_),
    .B_N(_06713_),
    .X(_07128_));
 sky130_fd_sc_hd__and4_2 _35177_ (.A(iX[49]),
    .B(iX[50]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_07129_));
 sky130_fd_sc_hd__a22oi_2 _35178_ (.A1(iX[50]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[49]),
    .Y(_07130_));
 sky130_fd_sc_hd__nor2_2 _35179_ (.A(_07129_),
    .B(_07130_),
    .Y(_07131_));
 sky130_fd_sc_hd__nand2_2 _35180_ (.A(iX[48]),
    .B(iY[61]),
    .Y(_07132_));
 sky130_fd_sc_hd__xnor2_2 _35181_ (.A(_07131_),
    .B(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__o21ba_2 _35182_ (.A1(_06710_),
    .A2(_06712_),
    .B1_N(_06709_),
    .X(_07134_));
 sky130_fd_sc_hd__xnor2_2 _35183_ (.A(_07133_),
    .B(_07134_),
    .Y(_07136_));
 sky130_fd_sc_hd__nand2_2 _35184_ (.A(iX[47]),
    .B(iY[62]),
    .Y(_07137_));
 sky130_fd_sc_hd__xor2_2 _35185_ (.A(_07136_),
    .B(_07137_),
    .X(_07138_));
 sky130_fd_sc_hd__a21oi_2 _35186_ (.A1(_07128_),
    .A2(_06718_),
    .B1(_07138_),
    .Y(_07139_));
 sky130_fd_sc_hd__and3_2 _35187_ (.A(_07128_),
    .B(_06718_),
    .C(_07138_),
    .X(_07140_));
 sky130_fd_sc_hd__nor2_2 _35188_ (.A(_07139_),
    .B(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__nand2_2 _35189_ (.A(iX[46]),
    .B(iY[63]),
    .Y(_07142_));
 sky130_fd_sc_hd__xnor2_2 _35190_ (.A(_07141_),
    .B(_07142_),
    .Y(_07143_));
 sky130_fd_sc_hd__or2b_2 _35191_ (.A(_06733_),
    .B_N(_06738_),
    .X(_07144_));
 sky130_fd_sc_hd__or2b_2 _35192_ (.A(_06732_),
    .B_N(_06739_),
    .X(_07145_));
 sky130_fd_sc_hd__and2b_2 _35193_ (.A_N(_06676_),
    .B(_06674_),
    .X(_07147_));
 sky130_fd_sc_hd__o21ba_2 _35194_ (.A1(_06735_),
    .A2(_06737_),
    .B1_N(_06734_),
    .X(_07148_));
 sky130_fd_sc_hd__o21ba_2 _35195_ (.A1(_06666_),
    .A2(_06668_),
    .B1_N(_06665_),
    .X(_07149_));
 sky130_fd_sc_hd__and4_2 _35196_ (.A(iX[52]),
    .B(iX[53]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_07150_));
 sky130_fd_sc_hd__a22oi_2 _35197_ (.A1(iX[53]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[52]),
    .Y(_07151_));
 sky130_fd_sc_hd__nor2_2 _35198_ (.A(_07150_),
    .B(_07151_),
    .Y(_07152_));
 sky130_fd_sc_hd__nand2_2 _35199_ (.A(iX[51]),
    .B(iY[58]),
    .Y(_07153_));
 sky130_fd_sc_hd__xnor2_2 _35200_ (.A(_07152_),
    .B(_07153_),
    .Y(_07154_));
 sky130_fd_sc_hd__xnor2_2 _35201_ (.A(_07149_),
    .B(_07154_),
    .Y(_07155_));
 sky130_fd_sc_hd__xnor2_2 _35202_ (.A(_07148_),
    .B(_07155_),
    .Y(_07156_));
 sky130_fd_sc_hd__o21a_2 _35203_ (.A1(_07147_),
    .A2(_06678_),
    .B1(_07156_),
    .X(_07158_));
 sky130_fd_sc_hd__nor3_2 _35204_ (.A(_07147_),
    .B(_06678_),
    .C(_07156_),
    .Y(_07159_));
 sky130_fd_sc_hd__a211oi_2 _35205_ (.A1(_07144_),
    .A2(_07145_),
    .B1(_07158_),
    .C1(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__o211a_2 _35206_ (.A1(_07158_),
    .A2(_07159_),
    .B1(_07144_),
    .C1(_07145_),
    .X(_07161_));
 sky130_fd_sc_hd__nor2_2 _35207_ (.A(_06741_),
    .B(_06743_),
    .Y(_07162_));
 sky130_fd_sc_hd__or3_2 _35208_ (.A(_07160_),
    .B(_07161_),
    .C(_07162_),
    .X(_07163_));
 sky130_fd_sc_hd__o21ai_2 _35209_ (.A1(_07160_),
    .A2(_07161_),
    .B1(_07162_),
    .Y(_07164_));
 sky130_fd_sc_hd__nand3_2 _35210_ (.A(_07143_),
    .B(_07163_),
    .C(_07164_),
    .Y(_07165_));
 sky130_fd_sc_hd__a21o_2 _35211_ (.A1(_07163_),
    .A2(_07164_),
    .B1(_07143_),
    .X(_07166_));
 sky130_fd_sc_hd__and2_2 _35212_ (.A(_07165_),
    .B(_07166_),
    .X(_07167_));
 sky130_fd_sc_hd__o21ai_2 _35213_ (.A1(_06698_),
    .A2(_06700_),
    .B1(_07167_),
    .Y(_07169_));
 sky130_fd_sc_hd__or3_2 _35214_ (.A(_06698_),
    .B(_06700_),
    .C(_07167_),
    .X(_07170_));
 sky130_fd_sc_hd__o211ai_2 _35215_ (.A1(_07127_),
    .A2(_06748_),
    .B1(_07169_),
    .C1(_07170_),
    .Y(_07171_));
 sky130_fd_sc_hd__a211o_2 _35216_ (.A1(_07169_),
    .A2(_07170_),
    .B1(_07127_),
    .C1(_06748_),
    .X(_07172_));
 sky130_fd_sc_hd__and3_2 _35217_ (.A(_07126_),
    .B(_07171_),
    .C(_07172_),
    .X(_07173_));
 sky130_fd_sc_hd__a21oi_2 _35218_ (.A1(_07171_),
    .A2(_07172_),
    .B1(_07126_),
    .Y(_07174_));
 sky130_fd_sc_hd__a211oi_2 _35219_ (.A1(_06705_),
    .A2(_06755_),
    .B1(_07173_),
    .C1(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__o211a_2 _35220_ (.A1(_07173_),
    .A2(_07174_),
    .B1(_06705_),
    .C1(_06755_),
    .X(_07176_));
 sky130_fd_sc_hd__a211oi_2 _35221_ (.A1(_07082_),
    .A2(_06753_),
    .B1(_07175_),
    .C1(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__o211a_2 _35222_ (.A1(_07175_),
    .A2(_07176_),
    .B1(_07082_),
    .C1(_06753_),
    .X(_07178_));
 sky130_fd_sc_hd__nor2_2 _35223_ (.A(_07177_),
    .B(_07178_),
    .Y(_07180_));
 sky130_fd_sc_hd__o21a_2 _35224_ (.A1(_06758_),
    .A2(_07081_),
    .B1(_07180_),
    .X(_07181_));
 sky130_fd_sc_hd__nor3_2 _35225_ (.A(_06758_),
    .B(_07081_),
    .C(_07180_),
    .Y(_07182_));
 sky130_fd_sc_hd__inv_2 _35226_ (.A(_06720_),
    .Y(_07183_));
 sky130_fd_sc_hd__a21oi_2 _35227_ (.A1(_07183_),
    .A2(_06722_),
    .B1(_06726_),
    .Y(_07184_));
 sky130_fd_sc_hd__or3_2 _35228_ (.A(_07181_),
    .B(_07182_),
    .C(_07184_),
    .X(_07185_));
 sky130_fd_sc_hd__o21ai_2 _35229_ (.A1(_07181_),
    .A2(_07182_),
    .B1(_07184_),
    .Y(_07186_));
 sky130_fd_sc_hd__nand2_2 _35230_ (.A(_07185_),
    .B(_07186_),
    .Y(_07187_));
 sky130_fd_sc_hd__o21a_2 _35231_ (.A1(_06636_),
    .A2(_06638_),
    .B1(_06763_),
    .X(_07188_));
 sky130_fd_sc_hd__a21oi_2 _35232_ (.A1(_06765_),
    .A2(_06766_),
    .B1(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__and2_2 _35233_ (.A(_07187_),
    .B(_07189_),
    .X(_07191_));
 sky130_fd_sc_hd__nor2_2 _35234_ (.A(_07187_),
    .B(_07189_),
    .Y(_07192_));
 sky130_fd_sc_hd__nor2_2 _35235_ (.A(_07191_),
    .B(_07192_),
    .Y(_07193_));
 sky130_fd_sc_hd__o21ba_2 _35236_ (.A1(_06770_),
    .A2(_06779_),
    .B1_N(_06769_),
    .X(_07194_));
 sky130_fd_sc_hd__xnor2_2 _35237_ (.A(_07193_),
    .B(_07194_),
    .Y(_07195_));
 sky130_fd_sc_hd__and3_2 _35238_ (.A(_07078_),
    .B(_07079_),
    .C(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__a21o_2 _35239_ (.A1(_07078_),
    .A2(_07079_),
    .B1(_07195_),
    .X(_07197_));
 sky130_fd_sc_hd__and2b_2 _35240_ (.A_N(_07196_),
    .B(_07197_),
    .X(_07198_));
 sky130_fd_sc_hd__xor2_2 _35241_ (.A(_14815_),
    .B(_07198_),
    .X(_07199_));
 sky130_fd_sc_hd__a21o_2 _35242_ (.A1(_14335_),
    .A2(_06921_),
    .B1(_06919_),
    .X(_07200_));
 sky130_fd_sc_hd__xor2_2 _35243_ (.A(_07199_),
    .B(_07200_),
    .X(_07202_));
 sky130_fd_sc_hd__a21oi_2 _35244_ (.A1(_06940_),
    .A2(_06931_),
    .B1(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__a31o_2 _35245_ (.A1(_06940_),
    .A2(_06931_),
    .A3(_07202_),
    .B1(_07203_),
    .X(_07204_));
 sky130_fd_sc_hd__nor2_2 _35246_ (.A(_14586_),
    .B(_07204_),
    .Y(_07205_));
 sky130_fd_sc_hd__nand2_2 _35247_ (.A(_14586_),
    .B(_07204_),
    .Y(_07206_));
 sky130_fd_sc_hd__and2b_2 _35248_ (.A_N(_07205_),
    .B(_07206_),
    .X(_07207_));
 sky130_fd_sc_hd__and2b_2 _35249_ (.A_N(_06939_),
    .B(_06936_),
    .X(_07208_));
 sky130_fd_sc_hd__nor2_2 _35250_ (.A(_06934_),
    .B(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__xnor2_2 _35251_ (.A(_07207_),
    .B(_07209_),
    .Y(oO[77]));
 sky130_fd_sc_hd__a31o_2 _35252_ (.A1(_06785_),
    .A2(_06789_),
    .A3(_06949_),
    .B1(_06947_),
    .X(_07210_));
 sky130_fd_sc_hd__or2_2 _35253_ (.A(_01034_),
    .B(_06399_),
    .X(_07212_));
 sky130_fd_sc_hd__a2bb2o_2 _35254_ (.A1_N(_02471_),
    .A2_N(_06786_),
    .B1(_04005_),
    .B2(_01033_),
    .X(_07213_));
 sky130_fd_sc_hd__nand2_2 _35255_ (.A(_07212_),
    .B(_07213_),
    .Y(_07214_));
 sky130_fd_sc_hd__xor2_2 _35256_ (.A(_07210_),
    .B(_07214_),
    .X(_07215_));
 sky130_fd_sc_hd__o22a_2 _35257_ (.A1(_05521_),
    .A2(_06797_),
    .B1(_05550_),
    .B2(_15155_),
    .X(_07216_));
 sky130_fd_sc_hd__and3b_2 _35258_ (.A_N(_05521_),
    .B(_03454_),
    .C(_06798_),
    .X(_07217_));
 sky130_fd_sc_hd__nor2_2 _35259_ (.A(_07216_),
    .B(_07217_),
    .Y(_07218_));
 sky130_fd_sc_hd__a21oi_2 _35260_ (.A1(_06957_),
    .A2(_06958_),
    .B1(_06955_),
    .Y(_07219_));
 sky130_fd_sc_hd__xnor2_2 _35261_ (.A(_07218_),
    .B(_07219_),
    .Y(_07220_));
 sky130_fd_sc_hd__xor2_2 _35262_ (.A(_06963_),
    .B(_07220_),
    .X(_07221_));
 sky130_fd_sc_hd__or4_2 _35263_ (.A(_05980_),
    .B(_05978_),
    .C(_04162_),
    .D(_05227_),
    .X(_07223_));
 sky130_fd_sc_hd__a22o_2 _35264_ (.A1(_06411_),
    .A2(_06822_),
    .B1(_06983_),
    .B2(_06414_),
    .X(_07224_));
 sky130_fd_sc_hd__nand2_2 _35265_ (.A(_07223_),
    .B(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__nand2_2 _35266_ (.A(_06813_),
    .B(_04138_),
    .Y(_07226_));
 sky130_fd_sc_hd__xnor2_2 _35267_ (.A(_07225_),
    .B(_07226_),
    .Y(_07227_));
 sky130_fd_sc_hd__nor2_2 _35268_ (.A(_01804_),
    .B(_05231_),
    .Y(_07228_));
 sky130_fd_sc_hd__xnor2_2 _35269_ (.A(_06978_),
    .B(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__nor2_2 _35270_ (.A(_04847_),
    .B(_05543_),
    .Y(_07230_));
 sky130_fd_sc_hd__xnor2_2 _35271_ (.A(_07229_),
    .B(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__o21a_2 _35272_ (.A1(_06982_),
    .A2(_06984_),
    .B1(_06979_),
    .X(_07232_));
 sky130_fd_sc_hd__or2_2 _35273_ (.A(_07231_),
    .B(_07232_),
    .X(_07234_));
 sky130_fd_sc_hd__nand2_2 _35274_ (.A(_07231_),
    .B(_07232_),
    .Y(_07235_));
 sky130_fd_sc_hd__nand2_2 _35275_ (.A(_07234_),
    .B(_07235_),
    .Y(_07236_));
 sky130_fd_sc_hd__xor2_2 _35276_ (.A(_07227_),
    .B(_07236_),
    .X(_07237_));
 sky130_fd_sc_hd__and2_2 _35277_ (.A(_07221_),
    .B(_07237_),
    .X(_07238_));
 sky130_fd_sc_hd__nor2_2 _35278_ (.A(_07221_),
    .B(_07237_),
    .Y(_07239_));
 sky130_fd_sc_hd__or2_2 _35279_ (.A(_07238_),
    .B(_07239_),
    .X(_07240_));
 sky130_fd_sc_hd__a21oi_2 _35280_ (.A1(_06969_),
    .A2(_06990_),
    .B1(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__and3_2 _35281_ (.A(_06969_),
    .B(_06990_),
    .C(_07240_),
    .X(_07242_));
 sky130_fd_sc_hd__or2_2 _35282_ (.A(_07241_),
    .B(_07242_),
    .X(_07243_));
 sky130_fd_sc_hd__inv_2 _35283_ (.A(_07243_),
    .Y(_07245_));
 sky130_fd_sc_hd__xnor2_2 _35284_ (.A(_07215_),
    .B(_07245_),
    .Y(_07246_));
 sky130_fd_sc_hd__a21boi_2 _35285_ (.A1(_06954_),
    .A2(_06997_),
    .B1_N(_06953_),
    .Y(_07247_));
 sky130_fd_sc_hd__xnor2_2 _35286_ (.A(_07246_),
    .B(_07247_),
    .Y(_07248_));
 sky130_fd_sc_hd__o21bai_2 _35287_ (.A1(_07029_),
    .A2(_07051_),
    .B1_N(_07050_),
    .Y(_07249_));
 sky130_fd_sc_hd__a21bo_2 _35288_ (.A1(_07011_),
    .A2(_07013_),
    .B1_N(_07010_),
    .X(_07250_));
 sky130_fd_sc_hd__or3_2 _35289_ (.A(_03389_),
    .B(_05931_),
    .C(_07009_),
    .X(_07251_));
 sky130_fd_sc_hd__buf_1 _35290_ (.A(_05931_),
    .X(_07252_));
 sky130_fd_sc_hd__a2bb2o_2 _35291_ (.A1_N(_01832_),
    .A2_N(_07252_),
    .B1(_04781_),
    .B2(_01040_),
    .X(_07253_));
 sky130_fd_sc_hd__nand2_2 _35292_ (.A(_07251_),
    .B(_07253_),
    .Y(_07254_));
 sky130_fd_sc_hd__nor2_2 _35293_ (.A(_03378_),
    .B(_05440_),
    .Y(_07256_));
 sky130_fd_sc_hd__xnor2_2 _35294_ (.A(_07254_),
    .B(_07256_),
    .Y(_07257_));
 sky130_fd_sc_hd__nand2_2 _35295_ (.A(_03024_),
    .B(_00567_),
    .Y(_07258_));
 sky130_fd_sc_hd__buf_1 _35296_ (.A(_02940_),
    .X(_07259_));
 sky130_fd_sc_hd__o22a_2 _35297_ (.A1(_04501_),
    .A2(_07259_),
    .B1(_02311_),
    .B2(_05983_),
    .X(_07260_));
 sky130_fd_sc_hd__o21bai_2 _35298_ (.A1(_07016_),
    .A2(_07258_),
    .B1_N(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__nand2_2 _35299_ (.A(_04837_),
    .B(_03327_),
    .Y(_07262_));
 sky130_fd_sc_hd__xnor2_2 _35300_ (.A(_07261_),
    .B(_07262_),
    .Y(_07263_));
 sky130_fd_sc_hd__o21a_2 _35301_ (.A1(_06853_),
    .A2(_07016_),
    .B1(_07018_),
    .X(_07264_));
 sky130_fd_sc_hd__nor2_2 _35302_ (.A(_07263_),
    .B(_07264_),
    .Y(_07265_));
 sky130_fd_sc_hd__and2_2 _35303_ (.A(_07263_),
    .B(_07264_),
    .X(_07267_));
 sky130_fd_sc_hd__nor2_2 _35304_ (.A(_07265_),
    .B(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__xnor2_2 _35305_ (.A(_07257_),
    .B(_07268_),
    .Y(_07269_));
 sky130_fd_sc_hd__a21o_2 _35306_ (.A1(_07015_),
    .A2(_07023_),
    .B1(_07022_),
    .X(_07270_));
 sky130_fd_sc_hd__xnor2_2 _35307_ (.A(_07269_),
    .B(_07270_),
    .Y(_07271_));
 sky130_fd_sc_hd__xnor2_2 _35308_ (.A(_07250_),
    .B(_07271_),
    .Y(_07272_));
 sky130_fd_sc_hd__and2b_2 _35309_ (.A_N(_07046_),
    .B(_07034_),
    .X(_07273_));
 sky130_fd_sc_hd__and2_2 _35310_ (.A(_07033_),
    .B(_07048_),
    .X(_07274_));
 sky130_fd_sc_hd__or2b_2 _35311_ (.A(_07044_),
    .B_N(_07038_),
    .X(_07275_));
 sky130_fd_sc_hd__a21bo_2 _35312_ (.A1(_07035_),
    .A2(_07045_),
    .B1_N(_07275_),
    .X(_07276_));
 sky130_fd_sc_hd__o21a_2 _35313_ (.A1(_06977_),
    .A2(_06988_),
    .B1(_06986_),
    .X(_07278_));
 sky130_fd_sc_hd__buf_1 _35314_ (.A(_06484_),
    .X(_07279_));
 sky130_fd_sc_hd__a31o_2 _35315_ (.A1(_03024_),
    .A2(_07279_),
    .A3(_07042_),
    .B1(_07040_),
    .X(_07280_));
 sky130_fd_sc_hd__nand2_2 _35316_ (.A(_06973_),
    .B(_06976_),
    .Y(_07281_));
 sky130_fd_sc_hd__and4_2 _35317_ (.A(_03973_),
    .B(_07039_),
    .C(_00662_),
    .D(_06488_),
    .X(_07282_));
 sky130_fd_sc_hd__a22o_2 _35318_ (.A1(_07039_),
    .A2(_06413_),
    .B1(_06488_),
    .B2(_03973_),
    .X(_07283_));
 sky130_fd_sc_hd__and2b_2 _35319_ (.A_N(_07282_),
    .B(_07283_),
    .X(_07284_));
 sky130_fd_sc_hd__nand2_2 _35320_ (.A(_05507_),
    .B(_06484_),
    .Y(_07285_));
 sky130_fd_sc_hd__xor2_2 _35321_ (.A(_07284_),
    .B(_07285_),
    .X(_07286_));
 sky130_fd_sc_hd__xnor2_2 _35322_ (.A(_07281_),
    .B(_07286_),
    .Y(_07287_));
 sky130_fd_sc_hd__xnor2_2 _35323_ (.A(_07280_),
    .B(_07287_),
    .Y(_07289_));
 sky130_fd_sc_hd__xnor2_2 _35324_ (.A(_07278_),
    .B(_07289_),
    .Y(_07290_));
 sky130_fd_sc_hd__xnor2_2 _35325_ (.A(_07276_),
    .B(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__o21a_2 _35326_ (.A1(_07273_),
    .A2(_07274_),
    .B1(_07291_),
    .X(_07292_));
 sky130_fd_sc_hd__nor3_2 _35327_ (.A(_07273_),
    .B(_07274_),
    .C(_07291_),
    .Y(_07293_));
 sky130_fd_sc_hd__nor2_2 _35328_ (.A(_07292_),
    .B(_07293_),
    .Y(_07294_));
 sky130_fd_sc_hd__xnor2_2 _35329_ (.A(_07272_),
    .B(_07294_),
    .Y(_07295_));
 sky130_fd_sc_hd__xnor2_2 _35330_ (.A(_06995_),
    .B(_07295_),
    .Y(_07296_));
 sky130_fd_sc_hd__xor2_2 _35331_ (.A(_07249_),
    .B(_07296_),
    .X(_07297_));
 sky130_fd_sc_hd__xor2_2 _35332_ (.A(_07248_),
    .B(_07297_),
    .X(_07298_));
 sky130_fd_sc_hd__a21boi_2 _35333_ (.A1(_07001_),
    .A2(_07055_),
    .B1_N(_07000_),
    .Y(_07300_));
 sky130_fd_sc_hd__xnor2_2 _35334_ (.A(_07298_),
    .B(_07300_),
    .Y(_07301_));
 sky130_fd_sc_hd__and2b_2 _35335_ (.A_N(_07054_),
    .B(_07005_),
    .X(_07302_));
 sky130_fd_sc_hd__a21o_2 _35336_ (.A1(_07006_),
    .A2(_07053_),
    .B1(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__and2b_2 _35337_ (.A_N(_07026_),
    .B(_07027_),
    .X(_07304_));
 sky130_fd_sc_hd__and2_2 _35338_ (.A(_07008_),
    .B(_07028_),
    .X(_07305_));
 sky130_fd_sc_hd__nor2_2 _35339_ (.A(_07304_),
    .B(_07305_),
    .Y(_07306_));
 sky130_fd_sc_hd__xnor2_2 _35340_ (.A(_07303_),
    .B(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__xnor2_2 _35341_ (.A(_07301_),
    .B(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__a21bo_2 _35342_ (.A1(_07060_),
    .A2(_07067_),
    .B1_N(_07059_),
    .X(_07309_));
 sky130_fd_sc_hd__xor2_2 _35343_ (.A(_07308_),
    .B(_07309_),
    .X(_07311_));
 sky130_fd_sc_hd__xnor2_2 _35344_ (.A(_07065_),
    .B(_07311_),
    .Y(_07312_));
 sky130_fd_sc_hd__a21boi_2 _35345_ (.A1(_06942_),
    .A2(_07072_),
    .B1_N(_07071_),
    .Y(_07313_));
 sky130_fd_sc_hd__xnor2_2 _35346_ (.A(_07312_),
    .B(_07313_),
    .Y(_07314_));
 sky130_fd_sc_hd__inv_2 _35347_ (.A(_07314_),
    .Y(_07315_));
 sky130_fd_sc_hd__or2b_2 _35348_ (.A(_06909_),
    .B_N(_07077_),
    .X(_07316_));
 sky130_fd_sc_hd__a21o_2 _35349_ (.A1(_06912_),
    .A2(_06915_),
    .B1(_07316_),
    .X(_07317_));
 sky130_fd_sc_hd__a21oi_2 _35350_ (.A1(_07075_),
    .A2(_07076_),
    .B1(_06907_),
    .Y(_07318_));
 sky130_fd_sc_hd__o21ba_2 _35351_ (.A1(_07075_),
    .A2(_07076_),
    .B1_N(_07318_),
    .X(_07319_));
 sky130_fd_sc_hd__nand2_2 _35352_ (.A(_07317_),
    .B(_07319_),
    .Y(_07320_));
 sky130_fd_sc_hd__xnor2_2 _35353_ (.A(_07315_),
    .B(_07320_),
    .Y(_07322_));
 sky130_fd_sc_hd__and2b_2 _35354_ (.A_N(_06702_),
    .B(_07125_),
    .X(_07323_));
 sky130_fd_sc_hd__or3_2 _35355_ (.A(_07083_),
    .B(_07121_),
    .C(_07122_),
    .X(_07324_));
 sky130_fd_sc_hd__and3_2 _35356_ (.A(iY[47]),
    .B(iX[63]),
    .C(_07086_),
    .X(_07325_));
 sky130_fd_sc_hd__a21o_2 _35357_ (.A1(iY[47]),
    .A2(iX[63]),
    .B1(_07086_),
    .X(_07326_));
 sky130_fd_sc_hd__and2b_2 _35358_ (.A_N(_07325_),
    .B(_07326_),
    .X(_07327_));
 sky130_fd_sc_hd__nand2_2 _35359_ (.A(iY[49]),
    .B(iX[61]),
    .Y(_07328_));
 sky130_fd_sc_hd__xnor2_2 _35360_ (.A(_07327_),
    .B(_07328_),
    .Y(_07329_));
 sky130_fd_sc_hd__o21ba_2 _35361_ (.A1(_07088_),
    .A2(_07090_),
    .B1_N(_07087_),
    .X(_07330_));
 sky130_fd_sc_hd__xnor2_2 _35362_ (.A(_07329_),
    .B(_07330_),
    .Y(_07331_));
 sky130_fd_sc_hd__o21a_2 _35363_ (.A1(_07093_),
    .A2(_07097_),
    .B1(_07331_),
    .X(_07333_));
 sky130_fd_sc_hd__nor3_2 _35364_ (.A(_07093_),
    .B(_07097_),
    .C(_07331_),
    .Y(_07334_));
 sky130_fd_sc_hd__nor2_2 _35365_ (.A(_07333_),
    .B(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__and4_2 _35366_ (.A(iY[53]),
    .B(iY[54]),
    .C(iX[56]),
    .D(iX[57]),
    .X(_07336_));
 sky130_fd_sc_hd__a22oi_2 _35367_ (.A1(iY[54]),
    .A2(iX[56]),
    .B1(iX[57]),
    .B2(iY[53]),
    .Y(_07337_));
 sky130_fd_sc_hd__nor2_2 _35368_ (.A(_07336_),
    .B(_07337_),
    .Y(_07338_));
 sky130_fd_sc_hd__nand2_2 _35369_ (.A(iX[55]),
    .B(iY[55]),
    .Y(_07339_));
 sky130_fd_sc_hd__xnor2_2 _35370_ (.A(_07338_),
    .B(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__and4_2 _35371_ (.A(iY[50]),
    .B(iY[51]),
    .C(iX[59]),
    .D(iX[60]),
    .X(_07341_));
 sky130_fd_sc_hd__a22oi_2 _35372_ (.A1(iY[51]),
    .A2(iX[59]),
    .B1(iX[60]),
    .B2(iY[50]),
    .Y(_07342_));
 sky130_fd_sc_hd__nor2_2 _35373_ (.A(_07341_),
    .B(_07342_),
    .Y(_07344_));
 sky130_fd_sc_hd__nand2_2 _35374_ (.A(iY[52]),
    .B(iX[58]),
    .Y(_07345_));
 sky130_fd_sc_hd__xnor2_2 _35375_ (.A(_07344_),
    .B(_07345_),
    .Y(_07346_));
 sky130_fd_sc_hd__o21ba_2 _35376_ (.A1(_07109_),
    .A2(_07111_),
    .B1_N(_07108_),
    .X(_07347_));
 sky130_fd_sc_hd__xnor2_2 _35377_ (.A(_07346_),
    .B(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__and2_2 _35378_ (.A(_07340_),
    .B(_07348_),
    .X(_07349_));
 sky130_fd_sc_hd__nor2_2 _35379_ (.A(_07340_),
    .B(_07348_),
    .Y(_07350_));
 sky130_fd_sc_hd__or2_2 _35380_ (.A(_07349_),
    .B(_07350_),
    .X(_07351_));
 sky130_fd_sc_hd__inv_2 _35381_ (.A(_07351_),
    .Y(_07352_));
 sky130_fd_sc_hd__xnor2_2 _35382_ (.A(_07335_),
    .B(_07352_),
    .Y(_07353_));
 sky130_fd_sc_hd__o21ba_2 _35383_ (.A1(_07100_),
    .A2(_07119_),
    .B1_N(_07353_),
    .X(_07355_));
 sky130_fd_sc_hd__or3b_2 _35384_ (.A(_07100_),
    .B(_07119_),
    .C_N(_07353_),
    .X(_07356_));
 sky130_fd_sc_hd__or2b_2 _35385_ (.A(_07355_),
    .B_N(_07356_),
    .X(_07357_));
 sky130_fd_sc_hd__xnor2_2 _35386_ (.A(_07324_),
    .B(_07357_),
    .Y(_07358_));
 sky130_fd_sc_hd__and4_2 _35387_ (.A(iX[50]),
    .B(iX[51]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_07359_));
 sky130_fd_sc_hd__a22oi_2 _35388_ (.A1(iX[51]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[50]),
    .Y(_07360_));
 sky130_fd_sc_hd__nor2_2 _35389_ (.A(_07359_),
    .B(_07360_),
    .Y(_07361_));
 sky130_fd_sc_hd__nand2_2 _35390_ (.A(iX[49]),
    .B(iY[61]),
    .Y(_07362_));
 sky130_fd_sc_hd__xnor2_2 _35391_ (.A(_07361_),
    .B(_07362_),
    .Y(_07363_));
 sky130_fd_sc_hd__o21ba_2 _35392_ (.A1(_07130_),
    .A2(_07132_),
    .B1_N(_07129_),
    .X(_07364_));
 sky130_fd_sc_hd__xnor2_2 _35393_ (.A(_07363_),
    .B(_07364_),
    .Y(_07366_));
 sky130_fd_sc_hd__and2_2 _35394_ (.A(iX[48]),
    .B(iY[62]),
    .X(_07367_));
 sky130_fd_sc_hd__or2_2 _35395_ (.A(_07366_),
    .B(_07367_),
    .X(_07368_));
 sky130_fd_sc_hd__nand2_2 _35396_ (.A(_07366_),
    .B(_07367_),
    .Y(_07369_));
 sky130_fd_sc_hd__and2b_2 _35397_ (.A_N(_07134_),
    .B(_07133_),
    .X(_07370_));
 sky130_fd_sc_hd__a31o_2 _35398_ (.A1(iX[47]),
    .A2(iY[62]),
    .A3(_07136_),
    .B1(_07370_),
    .X(_07371_));
 sky130_fd_sc_hd__nand3_2 _35399_ (.A(_07368_),
    .B(_07369_),
    .C(_07371_),
    .Y(_07372_));
 sky130_fd_sc_hd__a21o_2 _35400_ (.A1(_07368_),
    .A2(_07369_),
    .B1(_07371_),
    .X(_07373_));
 sky130_fd_sc_hd__nand2_2 _35401_ (.A(_07372_),
    .B(_07373_),
    .Y(_07374_));
 sky130_fd_sc_hd__nand2_2 _35402_ (.A(iX[47]),
    .B(iY[63]),
    .Y(_07375_));
 sky130_fd_sc_hd__nand2_2 _35403_ (.A(_07374_),
    .B(_07375_),
    .Y(_07377_));
 sky130_fd_sc_hd__or2_2 _35404_ (.A(_07374_),
    .B(_07375_),
    .X(_07378_));
 sky130_fd_sc_hd__and2_2 _35405_ (.A(_07377_),
    .B(_07378_),
    .X(_07379_));
 sky130_fd_sc_hd__or2b_2 _35406_ (.A(_07149_),
    .B_N(_07154_),
    .X(_07380_));
 sky130_fd_sc_hd__or2b_2 _35407_ (.A(_07148_),
    .B_N(_07155_),
    .X(_07381_));
 sky130_fd_sc_hd__and2b_2 _35408_ (.A_N(_07114_),
    .B(_07112_),
    .X(_07382_));
 sky130_fd_sc_hd__o21ba_2 _35409_ (.A1(_07151_),
    .A2(_07153_),
    .B1_N(_07150_),
    .X(_07383_));
 sky130_fd_sc_hd__o21ba_2 _35410_ (.A1(_07104_),
    .A2(_07106_),
    .B1_N(_07103_),
    .X(_07384_));
 sky130_fd_sc_hd__and4_2 _35411_ (.A(iX[53]),
    .B(iX[54]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_07385_));
 sky130_fd_sc_hd__a22oi_2 _35412_ (.A1(iX[54]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[53]),
    .Y(_07386_));
 sky130_fd_sc_hd__nor2_2 _35413_ (.A(_07385_),
    .B(_07386_),
    .Y(_07388_));
 sky130_fd_sc_hd__nand2_2 _35414_ (.A(iX[52]),
    .B(iY[58]),
    .Y(_07389_));
 sky130_fd_sc_hd__xnor2_2 _35415_ (.A(_07388_),
    .B(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__xnor2_2 _35416_ (.A(_07384_),
    .B(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__xnor2_2 _35417_ (.A(_07383_),
    .B(_07391_),
    .Y(_07392_));
 sky130_fd_sc_hd__o21a_2 _35418_ (.A1(_07382_),
    .A2(_07116_),
    .B1(_07392_),
    .X(_07393_));
 sky130_fd_sc_hd__nor3_2 _35419_ (.A(_07382_),
    .B(_07116_),
    .C(_07392_),
    .Y(_07394_));
 sky130_fd_sc_hd__a211oi_2 _35420_ (.A1(_07380_),
    .A2(_07381_),
    .B1(_07393_),
    .C1(_07394_),
    .Y(_07395_));
 sky130_fd_sc_hd__o211a_2 _35421_ (.A1(_07393_),
    .A2(_07394_),
    .B1(_07380_),
    .C1(_07381_),
    .X(_07396_));
 sky130_fd_sc_hd__nor2_2 _35422_ (.A(_07158_),
    .B(_07160_),
    .Y(_07397_));
 sky130_fd_sc_hd__or3_2 _35423_ (.A(_07395_),
    .B(_07396_),
    .C(_07397_),
    .X(_07399_));
 sky130_fd_sc_hd__o21ai_2 _35424_ (.A1(_07395_),
    .A2(_07396_),
    .B1(_07397_),
    .Y(_07400_));
 sky130_fd_sc_hd__nand3_2 _35425_ (.A(_07379_),
    .B(_07399_),
    .C(_07400_),
    .Y(_07401_));
 sky130_fd_sc_hd__a21o_2 _35426_ (.A1(_07399_),
    .A2(_07400_),
    .B1(_07379_),
    .X(_07402_));
 sky130_fd_sc_hd__and3_2 _35427_ (.A(_07121_),
    .B(_07401_),
    .C(_07402_),
    .X(_07403_));
 sky130_fd_sc_hd__a21oi_2 _35428_ (.A1(_07401_),
    .A2(_07402_),
    .B1(_07121_),
    .Y(_07404_));
 sky130_fd_sc_hd__a211oi_2 _35429_ (.A1(_07163_),
    .A2(_07165_),
    .B1(_07403_),
    .C1(_07404_),
    .Y(_07405_));
 sky130_fd_sc_hd__o211a_2 _35430_ (.A1(_07403_),
    .A2(_07404_),
    .B1(_07163_),
    .C1(_07165_),
    .X(_07406_));
 sky130_fd_sc_hd__or3_2 _35431_ (.A(_07358_),
    .B(_07405_),
    .C(_07406_),
    .X(_07407_));
 sky130_fd_sc_hd__o21ai_2 _35432_ (.A1(_07405_),
    .A2(_07406_),
    .B1(_07358_),
    .Y(_07408_));
 sky130_fd_sc_hd__o211a_2 _35433_ (.A1(_07323_),
    .A2(_07173_),
    .B1(_07407_),
    .C1(_07408_),
    .X(_07410_));
 sky130_fd_sc_hd__a211oi_2 _35434_ (.A1(_07407_),
    .A2(_07408_),
    .B1(_07323_),
    .C1(_07173_),
    .Y(_07411_));
 sky130_fd_sc_hd__or2_2 _35435_ (.A(_07410_),
    .B(_07411_),
    .X(_07412_));
 sky130_fd_sc_hd__nand2_2 _35436_ (.A(_07169_),
    .B(_07171_),
    .Y(_07413_));
 sky130_fd_sc_hd__xnor2_2 _35437_ (.A(_07412_),
    .B(_07413_),
    .Y(_07414_));
 sky130_fd_sc_hd__o21a_2 _35438_ (.A1(_07175_),
    .A2(_07177_),
    .B1(_07414_),
    .X(_07415_));
 sky130_fd_sc_hd__nor3_2 _35439_ (.A(_07175_),
    .B(_07177_),
    .C(_07414_),
    .Y(_07416_));
 sky130_fd_sc_hd__nor2_2 _35440_ (.A(_07415_),
    .B(_07416_),
    .Y(_07417_));
 sky130_fd_sc_hd__a31o_2 _35441_ (.A1(iX[46]),
    .A2(iY[63]),
    .A3(_07141_),
    .B1(_07139_),
    .X(_07418_));
 sky130_fd_sc_hd__xnor2_2 _35442_ (.A(_07417_),
    .B(_07418_),
    .Y(_07419_));
 sky130_fd_sc_hd__and2b_2 _35443_ (.A_N(_07181_),
    .B(_07185_),
    .X(_07421_));
 sky130_fd_sc_hd__nor2_2 _35444_ (.A(_07419_),
    .B(_07421_),
    .Y(_07422_));
 sky130_fd_sc_hd__and2_2 _35445_ (.A(_07419_),
    .B(_07421_),
    .X(_07423_));
 sky130_fd_sc_hd__nor2_2 _35446_ (.A(_07422_),
    .B(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__nand2_2 _35447_ (.A(_06771_),
    .B(_07193_),
    .Y(_07425_));
 sky130_fd_sc_hd__inv_2 _35448_ (.A(_07191_),
    .Y(_07426_));
 sky130_fd_sc_hd__a21oi_2 _35449_ (.A1(_06769_),
    .A2(_07426_),
    .B1(_07192_),
    .Y(_07427_));
 sky130_fd_sc_hd__o21ai_2 _35450_ (.A1(_06779_),
    .A2(_07425_),
    .B1(_07427_),
    .Y(_07428_));
 sky130_fd_sc_hd__xor2_2 _35451_ (.A(_07424_),
    .B(_07428_),
    .X(_07429_));
 sky130_fd_sc_hd__xor2_2 _35452_ (.A(_07322_),
    .B(_07429_),
    .X(_07430_));
 sky130_fd_sc_hd__xnor2_2 _35453_ (.A(_14925_),
    .B(_07430_),
    .Y(_07432_));
 sky130_fd_sc_hd__o21a_2 _35454_ (.A1(_14815_),
    .A2(_07196_),
    .B1(_07197_),
    .X(_07433_));
 sky130_fd_sc_hd__xnor2_2 _35455_ (.A(_07432_),
    .B(_07433_),
    .Y(_07434_));
 sky130_fd_sc_hd__or2b_2 _35456_ (.A(_07199_),
    .B_N(_07200_),
    .X(_07435_));
 sky130_fd_sc_hd__o31a_2 _35457_ (.A1(_06922_),
    .A2(_06924_),
    .A3(_07202_),
    .B1(_07435_),
    .X(_07436_));
 sky130_fd_sc_hd__o31a_2 _35458_ (.A1(_06925_),
    .A2(_06930_),
    .A3(_07202_),
    .B1(_07436_),
    .X(_07437_));
 sky130_fd_sc_hd__xor2_2 _35459_ (.A(_07434_),
    .B(_07437_),
    .X(_07438_));
 sky130_fd_sc_hd__nand2_2 _35460_ (.A(_15124_),
    .B(_07438_),
    .Y(_07439_));
 sky130_fd_sc_hd__or2_2 _35461_ (.A(_15124_),
    .B(_07438_),
    .X(_07440_));
 sky130_fd_sc_hd__nand2_2 _35462_ (.A(_07439_),
    .B(_07440_),
    .Y(_07441_));
 sky130_fd_sc_hd__a21o_2 _35463_ (.A1(_06934_),
    .A2(_07206_),
    .B1(_07205_),
    .X(_07443_));
 sky130_fd_sc_hd__a21oi_2 _35464_ (.A1(_07208_),
    .A2(_07207_),
    .B1(_07443_),
    .Y(_07444_));
 sky130_fd_sc_hd__xor2_2 _35465_ (.A(_07441_),
    .B(_07444_),
    .X(oO[78]));
 sky130_fd_sc_hd__or2_2 _35466_ (.A(_07432_),
    .B(_07433_),
    .X(_07445_));
 sky130_fd_sc_hd__o21ai_2 _35467_ (.A1(_07434_),
    .A2(_07437_),
    .B1(_07445_),
    .Y(_07446_));
 sky130_fd_sc_hd__or2_2 _35468_ (.A(_07312_),
    .B(_07313_),
    .X(_07447_));
 sky130_fd_sc_hd__a21o_2 _35469_ (.A1(_07317_),
    .A2(_07319_),
    .B1(_07314_),
    .X(_07448_));
 sky130_fd_sc_hd__o21a_2 _35470_ (.A1(_07304_),
    .A2(_07305_),
    .B1(_07303_),
    .X(_07449_));
 sky130_fd_sc_hd__and2b_2 _35471_ (.A_N(_07300_),
    .B(_07298_),
    .X(_07450_));
 sky130_fd_sc_hd__and2_2 _35472_ (.A(_07301_),
    .B(_07307_),
    .X(_07451_));
 sky130_fd_sc_hd__nor2_2 _35473_ (.A(_07246_),
    .B(_07247_),
    .Y(_07453_));
 sky130_fd_sc_hd__nor2_2 _35474_ (.A(_07248_),
    .B(_07297_),
    .Y(_07454_));
 sky130_fd_sc_hd__and2_2 _35475_ (.A(_07215_),
    .B(_07245_),
    .X(_07455_));
 sky130_fd_sc_hd__or2b_2 _35476_ (.A(_07219_),
    .B_N(_07218_),
    .X(_07456_));
 sky130_fd_sc_hd__nand2_2 _35477_ (.A(_15586_),
    .B(_03458_),
    .Y(_07457_));
 sky130_fd_sc_hd__and3b_2 _35478_ (.A_N(_05521_),
    .B(_04905_),
    .C(_07457_),
    .X(_07458_));
 sky130_fd_sc_hd__xnor2_2 _35479_ (.A(_07456_),
    .B(_07458_),
    .Y(_07459_));
 sky130_fd_sc_hd__or4_2 _35480_ (.A(_05980_),
    .B(_05978_),
    .C(_01070_),
    .D(_05543_),
    .X(_07460_));
 sky130_fd_sc_hd__buf_1 _35481_ (.A(_03438_),
    .X(_07461_));
 sky130_fd_sc_hd__a22o_2 _35482_ (.A1(_06411_),
    .A2(_02629_),
    .B1(_07461_),
    .B2(_06414_),
    .X(_07462_));
 sky130_fd_sc_hd__and2_2 _35483_ (.A(_07460_),
    .B(_07462_),
    .X(_07464_));
 sky130_fd_sc_hd__or3b_2 _35484_ (.A(_05500_),
    .B(_06816_),
    .C_N(_07464_),
    .X(_07465_));
 sky130_fd_sc_hd__a21o_2 _35485_ (.A1(_06813_),
    .A2(_06822_),
    .B1(_07464_),
    .X(_07466_));
 sky130_fd_sc_hd__nand2_2 _35486_ (.A(_07465_),
    .B(_07466_),
    .Y(_07467_));
 sky130_fd_sc_hd__or2_2 _35487_ (.A(_16606_),
    .B(_06797_),
    .X(_07468_));
 sky130_fd_sc_hd__or3_2 _35488_ (.A(_01804_),
    .B(_05231_),
    .C(_07468_),
    .X(_07469_));
 sky130_fd_sc_hd__a2bb2o_2 _35489_ (.A1_N(_16606_),
    .A2_N(_05231_),
    .B1(_03458_),
    .B2(_16934_),
    .X(_07470_));
 sky130_fd_sc_hd__nand2_2 _35490_ (.A(_07469_),
    .B(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__buf_1 _35491_ (.A(_02648_),
    .X(_07472_));
 sky130_fd_sc_hd__nand2_2 _35492_ (.A(_16614_),
    .B(_07472_),
    .Y(_07473_));
 sky130_fd_sc_hd__xnor2_2 _35493_ (.A(_07471_),
    .B(_07473_),
    .Y(_07475_));
 sky130_fd_sc_hd__nor2_2 _35494_ (.A(_16606_),
    .B(_06023_),
    .Y(_07476_));
 sky130_fd_sc_hd__a22o_2 _35495_ (.A1(_07476_),
    .A2(_07228_),
    .B1(_07229_),
    .B2(_07230_),
    .X(_07477_));
 sky130_fd_sc_hd__or2b_2 _35496_ (.A(_07475_),
    .B_N(_07477_),
    .X(_07478_));
 sky130_fd_sc_hd__or2b_2 _35497_ (.A(_07477_),
    .B_N(_07475_),
    .X(_07479_));
 sky130_fd_sc_hd__nand2_2 _35498_ (.A(_07478_),
    .B(_07479_),
    .Y(_07480_));
 sky130_fd_sc_hd__or2_2 _35499_ (.A(_07467_),
    .B(_07480_),
    .X(_07481_));
 sky130_fd_sc_hd__nand2_2 _35500_ (.A(_07467_),
    .B(_07480_),
    .Y(_07482_));
 sky130_fd_sc_hd__and2_2 _35501_ (.A(_07481_),
    .B(_07482_),
    .X(_07483_));
 sky130_fd_sc_hd__xnor2_2 _35502_ (.A(_07459_),
    .B(_07483_),
    .Y(_07484_));
 sky130_fd_sc_hd__a21oi_2 _35503_ (.A1(_06963_),
    .A2(_07220_),
    .B1(_07238_),
    .Y(_07486_));
 sky130_fd_sc_hd__nor2_2 _35504_ (.A(_07484_),
    .B(_07486_),
    .Y(_07487_));
 sky130_fd_sc_hd__and2_2 _35505_ (.A(_07484_),
    .B(_07486_),
    .X(_07488_));
 sky130_fd_sc_hd__nor2_2 _35506_ (.A(_07487_),
    .B(_07488_),
    .Y(_07489_));
 sky130_fd_sc_hd__a311o_2 _35507_ (.A1(_06785_),
    .A2(_06789_),
    .A3(_06949_),
    .B1(_07214_),
    .C1(_06947_),
    .X(_07490_));
 sky130_fd_sc_hd__or2_2 _35508_ (.A(_01808_),
    .B(_06399_),
    .X(_07491_));
 sky130_fd_sc_hd__o22a_2 _35509_ (.A1(_03378_),
    .A2(_06786_),
    .B1(_04901_),
    .B2(_15155_),
    .X(_07492_));
 sky130_fd_sc_hd__inv_2 _35510_ (.A(_07492_),
    .Y(_07493_));
 sky130_fd_sc_hd__nand2_2 _35511_ (.A(_07491_),
    .B(_07493_),
    .Y(_07494_));
 sky130_fd_sc_hd__nand3_2 _35512_ (.A(_07212_),
    .B(_07490_),
    .C(_07494_),
    .Y(_07495_));
 sky130_fd_sc_hd__a21o_2 _35513_ (.A1(_07212_),
    .A2(_07490_),
    .B1(_07494_),
    .X(_07497_));
 sky130_fd_sc_hd__nand3_2 _35514_ (.A(_07489_),
    .B(_07495_),
    .C(_07497_),
    .Y(_07498_));
 sky130_fd_sc_hd__a21o_2 _35515_ (.A1(_07495_),
    .A2(_07497_),
    .B1(_07489_),
    .X(_07499_));
 sky130_fd_sc_hd__nand3_2 _35516_ (.A(_07455_),
    .B(_07498_),
    .C(_07499_),
    .Y(_07500_));
 sky130_fd_sc_hd__a21o_2 _35517_ (.A1(_07498_),
    .A2(_07499_),
    .B1(_07455_),
    .X(_07501_));
 sky130_fd_sc_hd__o21bai_2 _35518_ (.A1(_07272_),
    .A2(_07293_),
    .B1_N(_07292_),
    .Y(_07502_));
 sky130_fd_sc_hd__o31a_2 _35519_ (.A1(_03378_),
    .A2(_05441_),
    .A3(_07254_),
    .B1(_07251_),
    .X(_07503_));
 sky130_fd_sc_hd__nand2_2 _35520_ (.A(_04837_),
    .B(_02928_),
    .Y(_07504_));
 sky130_fd_sc_hd__or3_2 _35521_ (.A(_03389_),
    .B(_07252_),
    .C(_07504_),
    .X(_07505_));
 sky130_fd_sc_hd__o21ai_2 _35522_ (.A1(_03389_),
    .A2(_07252_),
    .B1(_07504_),
    .Y(_07506_));
 sky130_fd_sc_hd__nand2_2 _35523_ (.A(_07505_),
    .B(_07506_),
    .Y(_07508_));
 sky130_fd_sc_hd__nor2_2 _35524_ (.A(_01832_),
    .B(_05440_),
    .Y(_07509_));
 sky130_fd_sc_hd__xnor2_2 _35525_ (.A(_07508_),
    .B(_07509_),
    .Y(_07510_));
 sky130_fd_sc_hd__nand2_2 _35526_ (.A(_05507_),
    .B(_05450_),
    .Y(_07511_));
 sky130_fd_sc_hd__xnor2_2 _35527_ (.A(_07258_),
    .B(_07511_),
    .Y(_07512_));
 sky130_fd_sc_hd__or3_2 _35528_ (.A(_05983_),
    .B(_00944_),
    .C(_07512_),
    .X(_07513_));
 sky130_fd_sc_hd__o21ai_2 _35529_ (.A1(_05983_),
    .A2(_00944_),
    .B1(_07512_),
    .Y(_07514_));
 sky130_fd_sc_hd__nand2_2 _35530_ (.A(_07513_),
    .B(_07514_),
    .Y(_07515_));
 sky130_fd_sc_hd__o22a_2 _35531_ (.A1(_07016_),
    .A2(_07258_),
    .B1(_07260_),
    .B2(_07262_),
    .X(_07516_));
 sky130_fd_sc_hd__nor2_2 _35532_ (.A(_07515_),
    .B(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__nand2_2 _35533_ (.A(_07515_),
    .B(_07516_),
    .Y(_07519_));
 sky130_fd_sc_hd__and2b_2 _35534_ (.A_N(_07517_),
    .B(_07519_),
    .X(_07520_));
 sky130_fd_sc_hd__xnor2_2 _35535_ (.A(_07510_),
    .B(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__a21o_2 _35536_ (.A1(_07257_),
    .A2(_07268_),
    .B1(_07265_),
    .X(_07522_));
 sky130_fd_sc_hd__xnor2_2 _35537_ (.A(_07521_),
    .B(_07522_),
    .Y(_07523_));
 sky130_fd_sc_hd__xnor2_2 _35538_ (.A(_07503_),
    .B(_07523_),
    .Y(_07524_));
 sky130_fd_sc_hd__nor2_2 _35539_ (.A(_07278_),
    .B(_07289_),
    .Y(_07525_));
 sky130_fd_sc_hd__and2b_2 _35540_ (.A_N(_07290_),
    .B(_07276_),
    .X(_07526_));
 sky130_fd_sc_hd__and2b_2 _35541_ (.A_N(_07286_),
    .B(_07281_),
    .X(_07527_));
 sky130_fd_sc_hd__a21o_2 _35542_ (.A1(_07280_),
    .A2(_07287_),
    .B1(_07527_),
    .X(_07528_));
 sky130_fd_sc_hd__o21ai_2 _35543_ (.A1(_07227_),
    .A2(_07236_),
    .B1(_07234_),
    .Y(_07530_));
 sky130_fd_sc_hd__a31o_2 _35544_ (.A1(_05507_),
    .A2(_06484_),
    .A3(_07283_),
    .B1(_07282_),
    .X(_07531_));
 sky130_fd_sc_hd__o21ai_2 _35545_ (.A1(_07225_),
    .A2(_07226_),
    .B1(_07223_),
    .Y(_07532_));
 sky130_fd_sc_hd__nand2_2 _35546_ (.A(_07039_),
    .B(_06413_),
    .Y(_07533_));
 sky130_fd_sc_hd__nand2_2 _35547_ (.A(_06488_),
    .B(_04138_),
    .Y(_07534_));
 sky130_fd_sc_hd__a22o_2 _35548_ (.A1(_06413_),
    .A2(_06488_),
    .B1(_04138_),
    .B2(_07039_),
    .X(_07535_));
 sky130_fd_sc_hd__o21ai_2 _35549_ (.A1(_07533_),
    .A2(_07534_),
    .B1(_07535_),
    .Y(_07536_));
 sky130_fd_sc_hd__nand2_2 _35550_ (.A(_03973_),
    .B(_06484_),
    .Y(_07537_));
 sky130_fd_sc_hd__xnor2_2 _35551_ (.A(_07536_),
    .B(_07537_),
    .Y(_07538_));
 sky130_fd_sc_hd__xnor2_2 _35552_ (.A(_07532_),
    .B(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__xnor2_2 _35553_ (.A(_07531_),
    .B(_07539_),
    .Y(_07541_));
 sky130_fd_sc_hd__xor2_2 _35554_ (.A(_07530_),
    .B(_07541_),
    .X(_07542_));
 sky130_fd_sc_hd__xnor2_2 _35555_ (.A(_07528_),
    .B(_07542_),
    .Y(_07543_));
 sky130_fd_sc_hd__o21a_2 _35556_ (.A1(_07525_),
    .A2(_07526_),
    .B1(_07543_),
    .X(_07544_));
 sky130_fd_sc_hd__nor3_2 _35557_ (.A(_07525_),
    .B(_07526_),
    .C(_07543_),
    .Y(_07545_));
 sky130_fd_sc_hd__nor2_2 _35558_ (.A(_07544_),
    .B(_07545_),
    .Y(_07546_));
 sky130_fd_sc_hd__xor2_2 _35559_ (.A(_07524_),
    .B(_07546_),
    .X(_07547_));
 sky130_fd_sc_hd__xnor2_2 _35560_ (.A(_07241_),
    .B(_07547_),
    .Y(_07548_));
 sky130_fd_sc_hd__xnor2_2 _35561_ (.A(_07502_),
    .B(_07548_),
    .Y(_07549_));
 sky130_fd_sc_hd__nand3_2 _35562_ (.A(_07500_),
    .B(_07501_),
    .C(_07549_),
    .Y(_07550_));
 sky130_fd_sc_hd__a21o_2 _35563_ (.A1(_07500_),
    .A2(_07501_),
    .B1(_07549_),
    .X(_07552_));
 sky130_fd_sc_hd__o211ai_2 _35564_ (.A1(_07453_),
    .A2(_07454_),
    .B1(_07550_),
    .C1(_07552_),
    .Y(_07553_));
 sky130_fd_sc_hd__a211o_2 _35565_ (.A1(_07550_),
    .A2(_07552_),
    .B1(_07453_),
    .C1(_07454_),
    .X(_07554_));
 sky130_fd_sc_hd__nand2_2 _35566_ (.A(_06995_),
    .B(_07295_),
    .Y(_07555_));
 sky130_fd_sc_hd__or2b_2 _35567_ (.A(_07296_),
    .B_N(_07249_),
    .X(_07556_));
 sky130_fd_sc_hd__and2b_2 _35568_ (.A_N(_07269_),
    .B(_07270_),
    .X(_07557_));
 sky130_fd_sc_hd__a21oi_2 _35569_ (.A1(_07250_),
    .A2(_07271_),
    .B1(_07557_),
    .Y(_07558_));
 sky130_fd_sc_hd__a21oi_2 _35570_ (.A1(_07555_),
    .A2(_07556_),
    .B1(_07558_),
    .Y(_07559_));
 sky130_fd_sc_hd__and3_2 _35571_ (.A(_07555_),
    .B(_07556_),
    .C(_07558_),
    .X(_07560_));
 sky130_fd_sc_hd__nor2_2 _35572_ (.A(_07559_),
    .B(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__nand3_2 _35573_ (.A(_07553_),
    .B(_07554_),
    .C(_07561_),
    .Y(_07563_));
 sky130_fd_sc_hd__a21o_2 _35574_ (.A1(_07553_),
    .A2(_07554_),
    .B1(_07561_),
    .X(_07564_));
 sky130_fd_sc_hd__o211ai_2 _35575_ (.A1(_07450_),
    .A2(_07451_),
    .B1(_07563_),
    .C1(_07564_),
    .Y(_07565_));
 sky130_fd_sc_hd__a211o_2 _35576_ (.A1(_07563_),
    .A2(_07564_),
    .B1(_07450_),
    .C1(_07451_),
    .X(_07566_));
 sky130_fd_sc_hd__and3_2 _35577_ (.A(_07449_),
    .B(_07565_),
    .C(_07566_),
    .X(_07567_));
 sky130_fd_sc_hd__a21oi_2 _35578_ (.A1(_07565_),
    .A2(_07566_),
    .B1(_07449_),
    .Y(_07568_));
 sky130_fd_sc_hd__or2b_2 _35579_ (.A(_07308_),
    .B_N(_07309_),
    .X(_07569_));
 sky130_fd_sc_hd__or2_2 _35580_ (.A(_07065_),
    .B(_07311_),
    .X(_07570_));
 sky130_fd_sc_hd__o211a_2 _35581_ (.A1(_07567_),
    .A2(_07568_),
    .B1(_07569_),
    .C1(_07570_),
    .X(_07571_));
 sky130_fd_sc_hd__a211o_2 _35582_ (.A1(_07569_),
    .A2(_07570_),
    .B1(_07567_),
    .C1(_07568_),
    .X(_07572_));
 sky130_fd_sc_hd__and2b_2 _35583_ (.A_N(_07571_),
    .B(_07572_),
    .X(_07574_));
 sky130_fd_sc_hd__nand3_2 _35584_ (.A(_07447_),
    .B(_07448_),
    .C(_07574_),
    .Y(_07575_));
 sky130_fd_sc_hd__a21o_4 _35585_ (.A1(_07447_),
    .A2(_07448_),
    .B1(_07574_),
    .X(_07576_));
 sky130_fd_sc_hd__and2_2 _35586_ (.A(_07417_),
    .B(_07418_),
    .X(_07577_));
 sky130_fd_sc_hd__and2b_2 _35587_ (.A_N(_07412_),
    .B(_07413_),
    .X(_07578_));
 sky130_fd_sc_hd__and2b_2 _35588_ (.A_N(_07330_),
    .B(_07329_),
    .X(_07579_));
 sky130_fd_sc_hd__nand2_2 _35589_ (.A(iY[48]),
    .B(iX[62]),
    .Y(_07580_));
 sky130_fd_sc_hd__nand2_2 _35590_ (.A(iY[49]),
    .B(iX[63]),
    .Y(_07581_));
 sky130_fd_sc_hd__a22o_2 _35591_ (.A1(iY[49]),
    .A2(iX[62]),
    .B1(iX[63]),
    .B2(iY[48]),
    .X(_07582_));
 sky130_fd_sc_hd__o21a_2 _35592_ (.A1(_07580_),
    .A2(_07581_),
    .B1(_07582_),
    .X(_07583_));
 sky130_fd_sc_hd__a31o_2 _35593_ (.A1(iY[49]),
    .A2(iX[61]),
    .A3(_07326_),
    .B1(_07325_),
    .X(_07585_));
 sky130_fd_sc_hd__nand2_2 _35594_ (.A(_07583_),
    .B(_07585_),
    .Y(_07586_));
 sky130_fd_sc_hd__or2_2 _35595_ (.A(_07583_),
    .B(_07585_),
    .X(_07587_));
 sky130_fd_sc_hd__and2_2 _35596_ (.A(_07586_),
    .B(_07587_),
    .X(_07588_));
 sky130_fd_sc_hd__or2_2 _35597_ (.A(_07579_),
    .B(_07588_),
    .X(_07589_));
 sky130_fd_sc_hd__nand2_2 _35598_ (.A(_07579_),
    .B(_07588_),
    .Y(_07590_));
 sky130_fd_sc_hd__nand2_2 _35599_ (.A(_07589_),
    .B(_07590_),
    .Y(_07591_));
 sky130_fd_sc_hd__and4_2 _35600_ (.A(iY[53]),
    .B(iY[54]),
    .C(iX[57]),
    .D(iX[58]),
    .X(_07592_));
 sky130_fd_sc_hd__a22oi_2 _35601_ (.A1(iY[54]),
    .A2(iX[57]),
    .B1(iX[58]),
    .B2(iY[53]),
    .Y(_07593_));
 sky130_fd_sc_hd__nor2_2 _35602_ (.A(_07592_),
    .B(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__nand2_2 _35603_ (.A(iY[55]),
    .B(iX[56]),
    .Y(_07596_));
 sky130_fd_sc_hd__xnor2_2 _35604_ (.A(_07594_),
    .B(_07596_),
    .Y(_07597_));
 sky130_fd_sc_hd__and4_2 _35605_ (.A(iY[50]),
    .B(iY[51]),
    .C(iX[60]),
    .D(iX[61]),
    .X(_07598_));
 sky130_fd_sc_hd__a22oi_2 _35606_ (.A1(iY[51]),
    .A2(iX[60]),
    .B1(iX[61]),
    .B2(iY[50]),
    .Y(_07599_));
 sky130_fd_sc_hd__nor2_2 _35607_ (.A(_07598_),
    .B(_07599_),
    .Y(_07600_));
 sky130_fd_sc_hd__nand2_2 _35608_ (.A(iY[52]),
    .B(iX[59]),
    .Y(_07601_));
 sky130_fd_sc_hd__xnor2_2 _35609_ (.A(_07600_),
    .B(_07601_),
    .Y(_07602_));
 sky130_fd_sc_hd__o21ba_2 _35610_ (.A1(_07342_),
    .A2(_07345_),
    .B1_N(_07341_),
    .X(_07603_));
 sky130_fd_sc_hd__xnor2_2 _35611_ (.A(_07602_),
    .B(_07603_),
    .Y(_07604_));
 sky130_fd_sc_hd__and2_2 _35612_ (.A(_07597_),
    .B(_07604_),
    .X(_07605_));
 sky130_fd_sc_hd__nor2_2 _35613_ (.A(_07597_),
    .B(_07604_),
    .Y(_07607_));
 sky130_fd_sc_hd__or2_2 _35614_ (.A(_07605_),
    .B(_07607_),
    .X(_07608_));
 sky130_fd_sc_hd__or2_2 _35615_ (.A(_07591_),
    .B(_07608_),
    .X(_07609_));
 sky130_fd_sc_hd__nand2_2 _35616_ (.A(_07591_),
    .B(_07608_),
    .Y(_07610_));
 sky130_fd_sc_hd__nand2_2 _35617_ (.A(_07609_),
    .B(_07610_),
    .Y(_07611_));
 sky130_fd_sc_hd__a21oi_2 _35618_ (.A1(_07335_),
    .A2(_07352_),
    .B1(_07333_),
    .Y(_07612_));
 sky130_fd_sc_hd__xnor2_2 _35619_ (.A(_07611_),
    .B(_07612_),
    .Y(_07613_));
 sky130_fd_sc_hd__or2b_2 _35620_ (.A(_07364_),
    .B_N(_07363_),
    .X(_07614_));
 sky130_fd_sc_hd__and4_2 _35621_ (.A(iX[51]),
    .B(iX[52]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_07615_));
 sky130_fd_sc_hd__a22oi_2 _35622_ (.A1(iX[52]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[51]),
    .Y(_07616_));
 sky130_fd_sc_hd__nor2_2 _35623_ (.A(_07615_),
    .B(_07616_),
    .Y(_07618_));
 sky130_fd_sc_hd__nand2_2 _35624_ (.A(iX[50]),
    .B(iY[61]),
    .Y(_07619_));
 sky130_fd_sc_hd__xnor2_2 _35625_ (.A(_07618_),
    .B(_07619_),
    .Y(_07620_));
 sky130_fd_sc_hd__o21ba_2 _35626_ (.A1(_07360_),
    .A2(_07362_),
    .B1_N(_07359_),
    .X(_07621_));
 sky130_fd_sc_hd__xnor2_2 _35627_ (.A(_07620_),
    .B(_07621_),
    .Y(_07622_));
 sky130_fd_sc_hd__nand2_2 _35628_ (.A(iX[49]),
    .B(iY[62]),
    .Y(_07623_));
 sky130_fd_sc_hd__xor2_2 _35629_ (.A(_07622_),
    .B(_07623_),
    .X(_07624_));
 sky130_fd_sc_hd__a21oi_2 _35630_ (.A1(_07614_),
    .A2(_07369_),
    .B1(_07624_),
    .Y(_07625_));
 sky130_fd_sc_hd__and3_2 _35631_ (.A(_07614_),
    .B(_07369_),
    .C(_07624_),
    .X(_07626_));
 sky130_fd_sc_hd__nor2_2 _35632_ (.A(_07625_),
    .B(_07626_),
    .Y(_07627_));
 sky130_fd_sc_hd__nand2_2 _35633_ (.A(iX[48]),
    .B(iY[63]),
    .Y(_07629_));
 sky130_fd_sc_hd__xnor2_2 _35634_ (.A(_07627_),
    .B(_07629_),
    .Y(_07630_));
 sky130_fd_sc_hd__or2b_2 _35635_ (.A(_07384_),
    .B_N(_07390_),
    .X(_07631_));
 sky130_fd_sc_hd__or2b_2 _35636_ (.A(_07383_),
    .B_N(_07391_),
    .X(_07632_));
 sky130_fd_sc_hd__and2b_2 _35637_ (.A_N(_07347_),
    .B(_07346_),
    .X(_07633_));
 sky130_fd_sc_hd__o21ba_2 _35638_ (.A1(_07386_),
    .A2(_07389_),
    .B1_N(_07385_),
    .X(_07634_));
 sky130_fd_sc_hd__o21ba_2 _35639_ (.A1(_07337_),
    .A2(_07339_),
    .B1_N(_07336_),
    .X(_07635_));
 sky130_fd_sc_hd__and4_2 _35640_ (.A(iX[54]),
    .B(iX[55]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_07636_));
 sky130_fd_sc_hd__a22oi_2 _35641_ (.A1(iX[55]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[54]),
    .Y(_07637_));
 sky130_fd_sc_hd__nor2_2 _35642_ (.A(_07636_),
    .B(_07637_),
    .Y(_07638_));
 sky130_fd_sc_hd__nand2_2 _35643_ (.A(iX[53]),
    .B(iY[58]),
    .Y(_07640_));
 sky130_fd_sc_hd__xnor2_2 _35644_ (.A(_07638_),
    .B(_07640_),
    .Y(_07641_));
 sky130_fd_sc_hd__xnor2_2 _35645_ (.A(_07635_),
    .B(_07641_),
    .Y(_07642_));
 sky130_fd_sc_hd__xnor2_2 _35646_ (.A(_07634_),
    .B(_07642_),
    .Y(_07643_));
 sky130_fd_sc_hd__o21a_2 _35647_ (.A1(_07633_),
    .A2(_07349_),
    .B1(_07643_),
    .X(_07644_));
 sky130_fd_sc_hd__nor3_2 _35648_ (.A(_07633_),
    .B(_07349_),
    .C(_07643_),
    .Y(_07645_));
 sky130_fd_sc_hd__a211oi_2 _35649_ (.A1(_07631_),
    .A2(_07632_),
    .B1(_07644_),
    .C1(_07645_),
    .Y(_07646_));
 sky130_fd_sc_hd__o211a_2 _35650_ (.A1(_07644_),
    .A2(_07645_),
    .B1(_07631_),
    .C1(_07632_),
    .X(_07647_));
 sky130_fd_sc_hd__nor2_2 _35651_ (.A(_07393_),
    .B(_07395_),
    .Y(_07648_));
 sky130_fd_sc_hd__or3_2 _35652_ (.A(_07646_),
    .B(_07647_),
    .C(_07648_),
    .X(_07649_));
 sky130_fd_sc_hd__o21ai_2 _35653_ (.A1(_07646_),
    .A2(_07647_),
    .B1(_07648_),
    .Y(_07651_));
 sky130_fd_sc_hd__nand3_2 _35654_ (.A(_07630_),
    .B(_07649_),
    .C(_07651_),
    .Y(_07652_));
 sky130_fd_sc_hd__a21o_2 _35655_ (.A1(_07649_),
    .A2(_07651_),
    .B1(_07630_),
    .X(_07653_));
 sky130_fd_sc_hd__and3_2 _35656_ (.A(_07355_),
    .B(_07652_),
    .C(_07653_),
    .X(_07654_));
 sky130_fd_sc_hd__a21oi_2 _35657_ (.A1(_07652_),
    .A2(_07653_),
    .B1(_07355_),
    .Y(_07655_));
 sky130_fd_sc_hd__a211oi_2 _35658_ (.A1(_07399_),
    .A2(_07401_),
    .B1(_07654_),
    .C1(_07655_),
    .Y(_07656_));
 sky130_fd_sc_hd__o211a_2 _35659_ (.A1(_07654_),
    .A2(_07655_),
    .B1(_07399_),
    .C1(_07401_),
    .X(_07657_));
 sky130_fd_sc_hd__or3_2 _35660_ (.A(_07613_),
    .B(_07656_),
    .C(_07657_),
    .X(_07658_));
 sky130_fd_sc_hd__o21ai_2 _35661_ (.A1(_07656_),
    .A2(_07657_),
    .B1(_07613_),
    .Y(_07659_));
 sky130_fd_sc_hd__o21ai_2 _35662_ (.A1(_07324_),
    .A2(_07357_),
    .B1(_07407_),
    .Y(_07660_));
 sky130_fd_sc_hd__nand3_2 _35663_ (.A(_07658_),
    .B(_07659_),
    .C(_07660_),
    .Y(_07662_));
 sky130_fd_sc_hd__a21o_2 _35664_ (.A1(_07658_),
    .A2(_07659_),
    .B1(_07660_),
    .X(_07663_));
 sky130_fd_sc_hd__o211ai_2 _35665_ (.A1(_07403_),
    .A2(_07405_),
    .B1(_07662_),
    .C1(_07663_),
    .Y(_07664_));
 sky130_fd_sc_hd__a211o_2 _35666_ (.A1(_07662_),
    .A2(_07663_),
    .B1(_07403_),
    .C1(_07405_),
    .X(_07665_));
 sky130_fd_sc_hd__o211a_2 _35667_ (.A1(_07410_),
    .A2(_07578_),
    .B1(_07664_),
    .C1(_07665_),
    .X(_07666_));
 sky130_fd_sc_hd__a211oi_2 _35668_ (.A1(_07664_),
    .A2(_07665_),
    .B1(_07410_),
    .C1(_07578_),
    .Y(_07667_));
 sky130_fd_sc_hd__a211oi_2 _35669_ (.A1(_07372_),
    .A2(_07378_),
    .B1(_07666_),
    .C1(_07667_),
    .Y(_07668_));
 sky130_fd_sc_hd__o211a_2 _35670_ (.A1(_07666_),
    .A2(_07667_),
    .B1(_07372_),
    .C1(_07378_),
    .X(_07669_));
 sky130_fd_sc_hd__nor2_2 _35671_ (.A(_07668_),
    .B(_07669_),
    .Y(_07670_));
 sky130_fd_sc_hd__or3_2 _35672_ (.A(_07415_),
    .B(_07577_),
    .C(_07670_),
    .X(_07671_));
 sky130_fd_sc_hd__o21ai_2 _35673_ (.A1(_07415_),
    .A2(_07577_),
    .B1(_07670_),
    .Y(_07673_));
 sky130_fd_sc_hd__and2_2 _35674_ (.A(_07671_),
    .B(_07673_),
    .X(_07674_));
 sky130_fd_sc_hd__a21oi_2 _35675_ (.A1(_07424_),
    .A2(_07428_),
    .B1(_07422_),
    .Y(_07675_));
 sky130_fd_sc_hd__xnor2_2 _35676_ (.A(_07674_),
    .B(_07675_),
    .Y(_07676_));
 sky130_fd_sc_hd__nand3_2 _35677_ (.A(_07575_),
    .B(_07576_),
    .C(_07676_),
    .Y(_07677_));
 sky130_fd_sc_hd__a21o_4 _35678_ (.A1(_07575_),
    .A2(_07576_),
    .B1(_07676_),
    .X(_07678_));
 sky130_fd_sc_hd__nand3_2 _35679_ (.A(_15460_),
    .B(_07677_),
    .C(_07678_),
    .Y(_07679_));
 sky130_fd_sc_hd__a21o_4 _35680_ (.A1(_07677_),
    .A2(_07678_),
    .B1(_15460_),
    .X(_07680_));
 sky130_fd_sc_hd__nor2_2 _35681_ (.A(_07322_),
    .B(_07429_),
    .Y(_07681_));
 sky130_fd_sc_hd__a21o_2 _35682_ (.A1(_14925_),
    .A2(_07430_),
    .B1(_07681_),
    .X(_07682_));
 sky130_fd_sc_hd__a21oi_2 _35683_ (.A1(_07679_),
    .A2(_07680_),
    .B1(_07682_),
    .Y(_07684_));
 sky130_fd_sc_hd__and3_4 _35684_ (.A(_07682_),
    .B(_07679_),
    .C(_07680_),
    .X(_07685_));
 sky130_fd_sc_hd__nor2_2 _35685_ (.A(_07684_),
    .B(_07685_),
    .Y(_07686_));
 sky130_fd_sc_hd__xnor2_2 _35686_ (.A(_07446_),
    .B(_07686_),
    .Y(_07687_));
 sky130_fd_sc_hd__xor2_2 _35687_ (.A(_15351_),
    .B(_07687_),
    .X(_07688_));
 sky130_fd_sc_hd__o21ai_2 _35688_ (.A1(_07441_),
    .A2(_07444_),
    .B1(_07439_),
    .Y(_07689_));
 sky130_fd_sc_hd__xnor2_2 _35689_ (.A(_07688_),
    .B(_07689_),
    .Y(oO[79]));
 sky130_fd_sc_hd__nand2_2 _35690_ (.A(_07315_),
    .B(_07574_),
    .Y(_07690_));
 sky130_fd_sc_hd__a211o_2 _35691_ (.A1(_06912_),
    .A2(_06915_),
    .B1(_07316_),
    .C1(_07690_),
    .X(_07691_));
 sky130_fd_sc_hd__or2_2 _35692_ (.A(_07447_),
    .B(_07571_),
    .X(_07692_));
 sky130_fd_sc_hd__o311a_2 _35693_ (.A1(_07314_),
    .A2(_07319_),
    .A3(_07571_),
    .B1(_07572_),
    .C1(_07692_),
    .X(_07694_));
 sky130_fd_sc_hd__inv_2 _35694_ (.A(_07500_),
    .Y(_07695_));
 sky130_fd_sc_hd__and3_2 _35695_ (.A(_07500_),
    .B(_07501_),
    .C(_07549_),
    .X(_07696_));
 sky130_fd_sc_hd__o22ai_2 _35696_ (.A1(_01832_),
    .A2(_06786_),
    .B1(_04901_),
    .B2(_05521_),
    .Y(_07697_));
 sky130_fd_sc_hd__o21ai_2 _35697_ (.A1(_02468_),
    .A2(_06399_),
    .B1(_07697_),
    .Y(_07698_));
 sky130_fd_sc_hd__a311o_2 _35698_ (.A1(_07212_),
    .A2(_07490_),
    .A3(_07491_),
    .B1(_07492_),
    .C1(_07698_),
    .X(_07699_));
 sky130_fd_sc_hd__o21a_2 _35699_ (.A1(_07212_),
    .A2(_07492_),
    .B1(_07491_),
    .X(_07700_));
 sky130_fd_sc_hd__o211ai_2 _35700_ (.A1(_07490_),
    .A2(_07492_),
    .B1(_07698_),
    .C1(_07700_),
    .Y(_07701_));
 sky130_fd_sc_hd__or4_2 _35701_ (.A(_05980_),
    .B(_17409_),
    .C(_05543_),
    .D(_04187_),
    .X(_07702_));
 sky130_fd_sc_hd__a22o_2 _35702_ (.A1(_06411_),
    .A2(_03438_),
    .B1(_02648_),
    .B2(_06414_),
    .X(_07703_));
 sky130_fd_sc_hd__and2_2 _35703_ (.A(_07702_),
    .B(_07703_),
    .X(_07705_));
 sky130_fd_sc_hd__or3b_2 _35704_ (.A(_05500_),
    .B(_05227_),
    .C_N(_07705_),
    .X(_07706_));
 sky130_fd_sc_hd__a21o_2 _35705_ (.A1(_06813_),
    .A2(_06983_),
    .B1(_07705_),
    .X(_07707_));
 sky130_fd_sc_hd__nand2_2 _35706_ (.A(_07706_),
    .B(_07707_),
    .Y(_07708_));
 sky130_fd_sc_hd__and3b_2 _35707_ (.A_N(_07468_),
    .B(_16934_),
    .C(_03454_),
    .X(_07709_));
 sky130_fd_sc_hd__o21a_2 _35708_ (.A1(_01804_),
    .A2(_05550_),
    .B1(_07468_),
    .X(_07710_));
 sky130_fd_sc_hd__nor2_2 _35709_ (.A(_07709_),
    .B(_07710_),
    .Y(_07711_));
 sky130_fd_sc_hd__nor2_2 _35710_ (.A(_04847_),
    .B(_05231_),
    .Y(_07712_));
 sky130_fd_sc_hd__xnor2_2 _35711_ (.A(_07711_),
    .B(_07712_),
    .Y(_07713_));
 sky130_fd_sc_hd__o21a_2 _35712_ (.A1(_07471_),
    .A2(_07473_),
    .B1(_07469_),
    .X(_07714_));
 sky130_fd_sc_hd__or2_2 _35713_ (.A(_07713_),
    .B(_07714_),
    .X(_07716_));
 sky130_fd_sc_hd__nand2_2 _35714_ (.A(_07713_),
    .B(_07714_),
    .Y(_07717_));
 sky130_fd_sc_hd__nand2_2 _35715_ (.A(_07716_),
    .B(_07717_),
    .Y(_07718_));
 sky130_fd_sc_hd__or2_2 _35716_ (.A(_07708_),
    .B(_07718_),
    .X(_07719_));
 sky130_fd_sc_hd__nand2_2 _35717_ (.A(_07708_),
    .B(_07718_),
    .Y(_07720_));
 sky130_fd_sc_hd__and2_2 _35718_ (.A(_07719_),
    .B(_07720_),
    .X(_07721_));
 sky130_fd_sc_hd__xnor2_2 _35719_ (.A(_07217_),
    .B(_07721_),
    .Y(_07722_));
 sky130_fd_sc_hd__and2b_2 _35720_ (.A_N(_07456_),
    .B(_07458_),
    .X(_07723_));
 sky130_fd_sc_hd__a31o_2 _35721_ (.A1(_07459_),
    .A2(_07481_),
    .A3(_07482_),
    .B1(_07723_),
    .X(_07724_));
 sky130_fd_sc_hd__xnor2_2 _35722_ (.A(_07722_),
    .B(_07724_),
    .Y(_07725_));
 sky130_fd_sc_hd__and3_2 _35723_ (.A(_07699_),
    .B(_07701_),
    .C(_07725_),
    .X(_07727_));
 sky130_fd_sc_hd__a21o_2 _35724_ (.A1(_07699_),
    .A2(_07701_),
    .B1(_07725_),
    .X(_07728_));
 sky130_fd_sc_hd__or3b_2 _35725_ (.A(_07498_),
    .B(_07727_),
    .C_N(_07728_),
    .X(_07729_));
 sky130_fd_sc_hd__nand3_2 _35726_ (.A(_07699_),
    .B(_07701_),
    .C(_07725_),
    .Y(_07730_));
 sky130_fd_sc_hd__a21bo_2 _35727_ (.A1(_07730_),
    .A2(_07728_),
    .B1_N(_07498_),
    .X(_07731_));
 sky130_fd_sc_hd__a21o_2 _35728_ (.A1(_07524_),
    .A2(_07546_),
    .B1(_07544_),
    .X(_07732_));
 sky130_fd_sc_hd__o31a_2 _35729_ (.A1(_01832_),
    .A2(_05441_),
    .A3(_07508_),
    .B1(_07505_),
    .X(_07733_));
 sky130_fd_sc_hd__or3_2 _35730_ (.A(_05983_),
    .B(_05931_),
    .C(_07504_),
    .X(_07734_));
 sky130_fd_sc_hd__a2bb2o_2 _35731_ (.A1_N(_04504_),
    .A2_N(_07252_),
    .B1(_04781_),
    .B2(_01837_),
    .X(_07735_));
 sky130_fd_sc_hd__nand2_2 _35732_ (.A(_07734_),
    .B(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__nor2_2 _35733_ (.A(_03389_),
    .B(_05440_),
    .Y(_07738_));
 sky130_fd_sc_hd__xnor2_2 _35734_ (.A(_07736_),
    .B(_07738_),
    .Y(_07739_));
 sky130_fd_sc_hd__nand2_2 _35735_ (.A(_03973_),
    .B(_00566_),
    .Y(_07740_));
 sky130_fd_sc_hd__o22a_2 _35736_ (.A1(_04862_),
    .A2(_07259_),
    .B1(_02311_),
    .B2(_05979_),
    .X(_07741_));
 sky130_fd_sc_hd__o21bai_2 _35737_ (.A1(_07511_),
    .A2(_07740_),
    .B1_N(_07741_),
    .Y(_07742_));
 sky130_fd_sc_hd__nand2_2 _35738_ (.A(_03024_),
    .B(_03327_),
    .Y(_07743_));
 sky130_fd_sc_hd__xnor2_2 _35739_ (.A(_07742_),
    .B(_07743_),
    .Y(_07744_));
 sky130_fd_sc_hd__o21a_2 _35740_ (.A1(_07258_),
    .A2(_07511_),
    .B1(_07513_),
    .X(_07745_));
 sky130_fd_sc_hd__nor2_2 _35741_ (.A(_07744_),
    .B(_07745_),
    .Y(_07746_));
 sky130_fd_sc_hd__and2_2 _35742_ (.A(_07744_),
    .B(_07745_),
    .X(_07747_));
 sky130_fd_sc_hd__nor2_2 _35743_ (.A(_07746_),
    .B(_07747_),
    .Y(_07749_));
 sky130_fd_sc_hd__xnor2_2 _35744_ (.A(_07739_),
    .B(_07749_),
    .Y(_07750_));
 sky130_fd_sc_hd__a21o_2 _35745_ (.A1(_07510_),
    .A2(_07519_),
    .B1(_07517_),
    .X(_07751_));
 sky130_fd_sc_hd__xnor2_2 _35746_ (.A(_07750_),
    .B(_07751_),
    .Y(_07752_));
 sky130_fd_sc_hd__xnor2_2 _35747_ (.A(_07733_),
    .B(_07752_),
    .Y(_07753_));
 sky130_fd_sc_hd__and2b_2 _35748_ (.A_N(_07538_),
    .B(_07532_),
    .X(_07754_));
 sky130_fd_sc_hd__and2_2 _35749_ (.A(_07531_),
    .B(_07539_),
    .X(_07755_));
 sky130_fd_sc_hd__nor2_2 _35750_ (.A(_07533_),
    .B(_07534_),
    .Y(_07756_));
 sky130_fd_sc_hd__a31o_2 _35751_ (.A1(_03973_),
    .A2(_07279_),
    .A3(_07535_),
    .B1(_07756_),
    .X(_07757_));
 sky130_fd_sc_hd__nand2_2 _35752_ (.A(_07460_),
    .B(_07465_),
    .Y(_07758_));
 sky130_fd_sc_hd__or3_2 _35753_ (.A(_06491_),
    .B(_06816_),
    .C(_07534_),
    .X(_07760_));
 sky130_fd_sc_hd__o21ai_2 _35754_ (.A1(_06491_),
    .A2(_06816_),
    .B1(_07534_),
    .Y(_07761_));
 sky130_fd_sc_hd__nand2_2 _35755_ (.A(_07760_),
    .B(_07761_),
    .Y(_07762_));
 sky130_fd_sc_hd__nand2_2 _35756_ (.A(_06413_),
    .B(_04469_),
    .Y(_07763_));
 sky130_fd_sc_hd__xnor2_2 _35757_ (.A(_07762_),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__xnor2_2 _35758_ (.A(_07758_),
    .B(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__xnor2_2 _35759_ (.A(_07757_),
    .B(_07765_),
    .Y(_07766_));
 sky130_fd_sc_hd__a21o_2 _35760_ (.A1(_07478_),
    .A2(_07481_),
    .B1(_07766_),
    .X(_07767_));
 sky130_fd_sc_hd__nand3_2 _35761_ (.A(_07478_),
    .B(_07481_),
    .C(_07766_),
    .Y(_07768_));
 sky130_fd_sc_hd__o211ai_2 _35762_ (.A1(_07754_),
    .A2(_07755_),
    .B1(_07767_),
    .C1(_07768_),
    .Y(_07769_));
 sky130_fd_sc_hd__a211o_2 _35763_ (.A1(_07767_),
    .A2(_07768_),
    .B1(_07754_),
    .C1(_07755_),
    .X(_07771_));
 sky130_fd_sc_hd__nand2_2 _35764_ (.A(_07769_),
    .B(_07771_),
    .Y(_07772_));
 sky130_fd_sc_hd__or2b_2 _35765_ (.A(_07541_),
    .B_N(_07530_),
    .X(_07773_));
 sky130_fd_sc_hd__or2b_2 _35766_ (.A(_07542_),
    .B_N(_07528_),
    .X(_07774_));
 sky130_fd_sc_hd__nand2_2 _35767_ (.A(_07773_),
    .B(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__xnor2_2 _35768_ (.A(_07772_),
    .B(_07775_),
    .Y(_07776_));
 sky130_fd_sc_hd__xnor2_2 _35769_ (.A(_07753_),
    .B(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__xnor2_2 _35770_ (.A(_07487_),
    .B(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__xor2_2 _35771_ (.A(_07732_),
    .B(_07778_),
    .X(_07779_));
 sky130_fd_sc_hd__nand3_2 _35772_ (.A(_07729_),
    .B(_07731_),
    .C(_07779_),
    .Y(_07780_));
 sky130_fd_sc_hd__a21o_2 _35773_ (.A1(_07729_),
    .A2(_07731_),
    .B1(_07779_),
    .X(_07782_));
 sky130_fd_sc_hd__o211a_2 _35774_ (.A1(_07695_),
    .A2(_07696_),
    .B1(_07780_),
    .C1(_07782_),
    .X(_07783_));
 sky130_fd_sc_hd__a211oi_2 _35775_ (.A1(_07780_),
    .A2(_07782_),
    .B1(_07695_),
    .C1(_07696_),
    .Y(_07784_));
 sky130_fd_sc_hd__nand2_2 _35776_ (.A(_07241_),
    .B(_07547_),
    .Y(_07785_));
 sky130_fd_sc_hd__or2b_2 _35777_ (.A(_07548_),
    .B_N(_07502_),
    .X(_07786_));
 sky130_fd_sc_hd__and2b_2 _35778_ (.A_N(_07521_),
    .B(_07522_),
    .X(_07787_));
 sky130_fd_sc_hd__and2b_2 _35779_ (.A_N(_07503_),
    .B(_07523_),
    .X(_07788_));
 sky130_fd_sc_hd__nor2_2 _35780_ (.A(_07787_),
    .B(_07788_),
    .Y(_07789_));
 sky130_fd_sc_hd__a21oi_2 _35781_ (.A1(_07785_),
    .A2(_07786_),
    .B1(_07789_),
    .Y(_07790_));
 sky130_fd_sc_hd__and3_2 _35782_ (.A(_07785_),
    .B(_07786_),
    .C(_07789_),
    .X(_07791_));
 sky130_fd_sc_hd__or2_2 _35783_ (.A(_07790_),
    .B(_07791_),
    .X(_07793_));
 sky130_fd_sc_hd__nor3_2 _35784_ (.A(_07783_),
    .B(_07784_),
    .C(_07793_),
    .Y(_07794_));
 sky130_fd_sc_hd__o21a_2 _35785_ (.A1(_07783_),
    .A2(_07784_),
    .B1(_07793_),
    .X(_07795_));
 sky130_fd_sc_hd__a211o_2 _35786_ (.A1(_07553_),
    .A2(_07563_),
    .B1(_07794_),
    .C1(_07795_),
    .X(_07796_));
 sky130_fd_sc_hd__o211ai_2 _35787_ (.A1(_07794_),
    .A2(_07795_),
    .B1(_07553_),
    .C1(_07563_),
    .Y(_07797_));
 sky130_fd_sc_hd__and2_2 _35788_ (.A(_07796_),
    .B(_07797_),
    .X(_07798_));
 sky130_fd_sc_hd__nand2_2 _35789_ (.A(_07559_),
    .B(_07798_),
    .Y(_07799_));
 sky130_fd_sc_hd__or2_2 _35790_ (.A(_07559_),
    .B(_07798_),
    .X(_07800_));
 sky130_fd_sc_hd__nand2_2 _35791_ (.A(_07799_),
    .B(_07800_),
    .Y(_07801_));
 sky130_fd_sc_hd__inv_2 _35792_ (.A(_07565_),
    .Y(_07802_));
 sky130_fd_sc_hd__nor2_2 _35793_ (.A(_07802_),
    .B(_07567_),
    .Y(_07804_));
 sky130_fd_sc_hd__or2_2 _35794_ (.A(_07801_),
    .B(_07804_),
    .X(_07805_));
 sky130_fd_sc_hd__nand2_2 _35795_ (.A(_07801_),
    .B(_07804_),
    .Y(_07806_));
 sky130_fd_sc_hd__nand2_2 _35796_ (.A(_07805_),
    .B(_07806_),
    .Y(_07807_));
 sky130_fd_sc_hd__a21oi_2 _35797_ (.A1(_07691_),
    .A2(_07694_),
    .B1(_07807_),
    .Y(_07808_));
 sky130_fd_sc_hd__and3_2 _35798_ (.A(_07807_),
    .B(_07691_),
    .C(_07694_),
    .X(_07809_));
 sky130_fd_sc_hd__nor2_2 _35799_ (.A(_07808_),
    .B(_07809_),
    .Y(_07810_));
 sky130_fd_sc_hd__o21ba_2 _35800_ (.A1(_07626_),
    .A2(_07629_),
    .B1_N(_07625_),
    .X(_07811_));
 sky130_fd_sc_hd__nor2_2 _35801_ (.A(_07086_),
    .B(_07581_),
    .Y(_07812_));
 sky130_fd_sc_hd__xor2_2 _35802_ (.A(_07586_),
    .B(_07812_),
    .X(_07813_));
 sky130_fd_sc_hd__and4_2 _35803_ (.A(iY[53]),
    .B(iY[54]),
    .C(iX[58]),
    .D(iX[59]),
    .X(_07815_));
 sky130_fd_sc_hd__a22oi_2 _35804_ (.A1(iY[54]),
    .A2(iX[58]),
    .B1(iX[59]),
    .B2(iY[53]),
    .Y(_07816_));
 sky130_fd_sc_hd__nor2_2 _35805_ (.A(_07815_),
    .B(_07816_),
    .Y(_07817_));
 sky130_fd_sc_hd__nand2_2 _35806_ (.A(iY[55]),
    .B(iX[57]),
    .Y(_07818_));
 sky130_fd_sc_hd__xnor2_2 _35807_ (.A(_07817_),
    .B(_07818_),
    .Y(_07819_));
 sky130_fd_sc_hd__and2_2 _35808_ (.A(iY[51]),
    .B(iX[62]),
    .X(_07820_));
 sky130_fd_sc_hd__and3_2 _35809_ (.A(iY[50]),
    .B(iX[61]),
    .C(_07820_),
    .X(_07821_));
 sky130_fd_sc_hd__a22oi_2 _35810_ (.A1(iY[51]),
    .A2(iX[61]),
    .B1(iX[62]),
    .B2(iY[50]),
    .Y(_07822_));
 sky130_fd_sc_hd__nand2_2 _35811_ (.A(iY[52]),
    .B(iX[60]),
    .Y(_07823_));
 sky130_fd_sc_hd__o21a_2 _35812_ (.A1(_07821_),
    .A2(_07822_),
    .B1(_07823_),
    .X(_07824_));
 sky130_fd_sc_hd__nor3_2 _35813_ (.A(_07821_),
    .B(_07822_),
    .C(_07823_),
    .Y(_07826_));
 sky130_fd_sc_hd__nor2_2 _35814_ (.A(_07824_),
    .B(_07826_),
    .Y(_07827_));
 sky130_fd_sc_hd__o21ba_2 _35815_ (.A1(_07599_),
    .A2(_07601_),
    .B1_N(_07598_),
    .X(_07828_));
 sky130_fd_sc_hd__xnor2_2 _35816_ (.A(_07827_),
    .B(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__and2_2 _35817_ (.A(_07819_),
    .B(_07829_),
    .X(_07830_));
 sky130_fd_sc_hd__nor2_2 _35818_ (.A(_07819_),
    .B(_07829_),
    .Y(_07831_));
 sky130_fd_sc_hd__or2_2 _35819_ (.A(_07830_),
    .B(_07831_),
    .X(_07832_));
 sky130_fd_sc_hd__nor2_2 _35820_ (.A(_07813_),
    .B(_07832_),
    .Y(_07833_));
 sky130_fd_sc_hd__and2_2 _35821_ (.A(_07813_),
    .B(_07832_),
    .X(_07834_));
 sky130_fd_sc_hd__a211o_2 _35822_ (.A1(_07590_),
    .A2(_07609_),
    .B1(_07833_),
    .C1(_07834_),
    .X(_07835_));
 sky130_fd_sc_hd__o211ai_2 _35823_ (.A1(_07833_),
    .A2(_07834_),
    .B1(_07590_),
    .C1(_07609_),
    .Y(_07837_));
 sky130_fd_sc_hd__nor2_2 _35824_ (.A(_07611_),
    .B(_07612_),
    .Y(_07838_));
 sky130_fd_sc_hd__and4_2 _35825_ (.A(iX[52]),
    .B(iX[53]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_07839_));
 sky130_fd_sc_hd__a22oi_2 _35826_ (.A1(iX[53]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[52]),
    .Y(_07840_));
 sky130_fd_sc_hd__nor2_2 _35827_ (.A(_07839_),
    .B(_07840_),
    .Y(_07841_));
 sky130_fd_sc_hd__nand2_2 _35828_ (.A(iX[51]),
    .B(iY[61]),
    .Y(_07842_));
 sky130_fd_sc_hd__xnor2_2 _35829_ (.A(_07841_),
    .B(_07842_),
    .Y(_07843_));
 sky130_fd_sc_hd__o21ba_2 _35830_ (.A1(_07616_),
    .A2(_07619_),
    .B1_N(_07615_),
    .X(_07844_));
 sky130_fd_sc_hd__xnor2_2 _35831_ (.A(_07843_),
    .B(_07844_),
    .Y(_07845_));
 sky130_fd_sc_hd__and2_2 _35832_ (.A(iX[50]),
    .B(iY[62]),
    .X(_07846_));
 sky130_fd_sc_hd__or2_2 _35833_ (.A(_07845_),
    .B(_07846_),
    .X(_07848_));
 sky130_fd_sc_hd__nand2_2 _35834_ (.A(_07845_),
    .B(_07846_),
    .Y(_07849_));
 sky130_fd_sc_hd__and2b_2 _35835_ (.A_N(_07621_),
    .B(_07620_),
    .X(_07850_));
 sky130_fd_sc_hd__a31o_2 _35836_ (.A1(iX[49]),
    .A2(iY[62]),
    .A3(_07622_),
    .B1(_07850_),
    .X(_07851_));
 sky130_fd_sc_hd__nand3_2 _35837_ (.A(_07848_),
    .B(_07849_),
    .C(_07851_),
    .Y(_07852_));
 sky130_fd_sc_hd__a21o_2 _35838_ (.A1(_07848_),
    .A2(_07849_),
    .B1(_07851_),
    .X(_07853_));
 sky130_fd_sc_hd__nand2_2 _35839_ (.A(_07852_),
    .B(_07853_),
    .Y(_07854_));
 sky130_fd_sc_hd__nand2_2 _35840_ (.A(iX[49]),
    .B(iY[63]),
    .Y(_07855_));
 sky130_fd_sc_hd__nand2_2 _35841_ (.A(_07854_),
    .B(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__or2_2 _35842_ (.A(_07854_),
    .B(_07855_),
    .X(_07857_));
 sky130_fd_sc_hd__and2_2 _35843_ (.A(_07856_),
    .B(_07857_),
    .X(_07859_));
 sky130_fd_sc_hd__or2b_2 _35844_ (.A(_07635_),
    .B_N(_07641_),
    .X(_07860_));
 sky130_fd_sc_hd__or2b_2 _35845_ (.A(_07634_),
    .B_N(_07642_),
    .X(_07861_));
 sky130_fd_sc_hd__and2b_2 _35846_ (.A_N(_07603_),
    .B(_07602_),
    .X(_07862_));
 sky130_fd_sc_hd__o21ba_2 _35847_ (.A1(_07637_),
    .A2(_07640_),
    .B1_N(_07636_),
    .X(_07863_));
 sky130_fd_sc_hd__o21ba_2 _35848_ (.A1(_07593_),
    .A2(_07596_),
    .B1_N(_07592_),
    .X(_07864_));
 sky130_fd_sc_hd__and4_2 _35849_ (.A(iX[55]),
    .B(iX[56]),
    .C(iY[56]),
    .D(iY[57]),
    .X(_07865_));
 sky130_fd_sc_hd__a22oi_2 _35850_ (.A1(iX[56]),
    .A2(iY[56]),
    .B1(iY[57]),
    .B2(iX[55]),
    .Y(_07866_));
 sky130_fd_sc_hd__nor2_2 _35851_ (.A(_07865_),
    .B(_07866_),
    .Y(_07867_));
 sky130_fd_sc_hd__nand2_2 _35852_ (.A(iX[54]),
    .B(iY[58]),
    .Y(_07868_));
 sky130_fd_sc_hd__xnor2_2 _35853_ (.A(_07867_),
    .B(_07868_),
    .Y(_07870_));
 sky130_fd_sc_hd__xnor2_2 _35854_ (.A(_07864_),
    .B(_07870_),
    .Y(_07871_));
 sky130_fd_sc_hd__xnor2_2 _35855_ (.A(_07863_),
    .B(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__o21a_2 _35856_ (.A1(_07862_),
    .A2(_07605_),
    .B1(_07872_),
    .X(_07873_));
 sky130_fd_sc_hd__nor3_2 _35857_ (.A(_07862_),
    .B(_07605_),
    .C(_07872_),
    .Y(_07874_));
 sky130_fd_sc_hd__a211oi_2 _35858_ (.A1(_07860_),
    .A2(_07861_),
    .B1(_07873_),
    .C1(_07874_),
    .Y(_07875_));
 sky130_fd_sc_hd__o211a_2 _35859_ (.A1(_07873_),
    .A2(_07874_),
    .B1(_07860_),
    .C1(_07861_),
    .X(_07876_));
 sky130_fd_sc_hd__nor2_2 _35860_ (.A(_07644_),
    .B(_07646_),
    .Y(_07877_));
 sky130_fd_sc_hd__or3_2 _35861_ (.A(_07875_),
    .B(_07876_),
    .C(_07877_),
    .X(_07878_));
 sky130_fd_sc_hd__o21ai_2 _35862_ (.A1(_07875_),
    .A2(_07876_),
    .B1(_07877_),
    .Y(_07879_));
 sky130_fd_sc_hd__nand3_2 _35863_ (.A(_07859_),
    .B(_07878_),
    .C(_07879_),
    .Y(_07881_));
 sky130_fd_sc_hd__a21o_2 _35864_ (.A1(_07878_),
    .A2(_07879_),
    .B1(_07859_),
    .X(_07882_));
 sky130_fd_sc_hd__nand3_2 _35865_ (.A(_07838_),
    .B(_07881_),
    .C(_07882_),
    .Y(_07883_));
 sky130_fd_sc_hd__a21o_2 _35866_ (.A1(_07881_),
    .A2(_07882_),
    .B1(_07838_),
    .X(_07884_));
 sky130_fd_sc_hd__nand2_2 _35867_ (.A(_07883_),
    .B(_07884_),
    .Y(_07885_));
 sky130_fd_sc_hd__a21o_2 _35868_ (.A1(_07649_),
    .A2(_07652_),
    .B1(_07885_),
    .X(_07886_));
 sky130_fd_sc_hd__nand3_2 _35869_ (.A(_07649_),
    .B(_07652_),
    .C(_07885_),
    .Y(_07887_));
 sky130_fd_sc_hd__and4_2 _35870_ (.A(_07835_),
    .B(_07837_),
    .C(_07886_),
    .D(_07887_),
    .X(_07888_));
 sky130_fd_sc_hd__a22oi_2 _35871_ (.A1(_07835_),
    .A2(_07837_),
    .B1(_07886_),
    .B2(_07887_),
    .Y(_07889_));
 sky130_fd_sc_hd__or3_2 _35872_ (.A(_07658_),
    .B(_07888_),
    .C(_07889_),
    .X(_07890_));
 sky130_fd_sc_hd__o21ai_2 _35873_ (.A1(_07888_),
    .A2(_07889_),
    .B1(_07658_),
    .Y(_07892_));
 sky130_fd_sc_hd__o211ai_2 _35874_ (.A1(_07654_),
    .A2(_07656_),
    .B1(_07890_),
    .C1(_07892_),
    .Y(_07893_));
 sky130_fd_sc_hd__a211o_2 _35875_ (.A1(_07890_),
    .A2(_07892_),
    .B1(_07654_),
    .C1(_07656_),
    .X(_07894_));
 sky130_fd_sc_hd__and2_2 _35876_ (.A(_07893_),
    .B(_07894_),
    .X(_07895_));
 sky130_fd_sc_hd__nand2_2 _35877_ (.A(_07662_),
    .B(_07664_),
    .Y(_07896_));
 sky130_fd_sc_hd__xor2_2 _35878_ (.A(_07895_),
    .B(_07896_),
    .X(_07897_));
 sky130_fd_sc_hd__and2b_2 _35879_ (.A_N(_07811_),
    .B(_07897_),
    .X(_07898_));
 sky130_fd_sc_hd__and2b_2 _35880_ (.A_N(_07897_),
    .B(_07811_),
    .X(_07899_));
 sky130_fd_sc_hd__or2_2 _35881_ (.A(_07898_),
    .B(_07899_),
    .X(_07900_));
 sky130_fd_sc_hd__nor2_2 _35882_ (.A(_07666_),
    .B(_07668_),
    .Y(_07901_));
 sky130_fd_sc_hd__nor2_2 _35883_ (.A(_07900_),
    .B(_07901_),
    .Y(_07903_));
 sky130_fd_sc_hd__and2_2 _35884_ (.A(_07900_),
    .B(_07901_),
    .X(_07904_));
 sky130_fd_sc_hd__or2_2 _35885_ (.A(_07903_),
    .B(_07904_),
    .X(_07905_));
 sky130_fd_sc_hd__nand2_2 _35886_ (.A(_07424_),
    .B(_07674_),
    .Y(_07906_));
 sky130_fd_sc_hd__a211o_2 _35887_ (.A1(_06774_),
    .A2(_06778_),
    .B1(_07425_),
    .C1(_07906_),
    .X(_07907_));
 sky130_fd_sc_hd__nand2_2 _35888_ (.A(_07422_),
    .B(_07671_),
    .Y(_07908_));
 sky130_fd_sc_hd__o211a_2 _35889_ (.A1(_07427_),
    .A2(_07906_),
    .B1(_07908_),
    .C1(_07673_),
    .X(_07909_));
 sky130_fd_sc_hd__and2_2 _35890_ (.A(_07907_),
    .B(_07909_),
    .X(_07910_));
 sky130_fd_sc_hd__xor2_2 _35891_ (.A(_07905_),
    .B(_07910_),
    .X(_07911_));
 sky130_fd_sc_hd__xnor2_2 _35892_ (.A(_07810_),
    .B(_07911_),
    .Y(_07912_));
 sky130_fd_sc_hd__xor2_2 _35893_ (.A(_15575_),
    .B(_07912_),
    .X(_07914_));
 sky130_fd_sc_hd__a21boi_2 _35894_ (.A1(_15460_),
    .A2(_07677_),
    .B1_N(_07678_),
    .Y(_07915_));
 sky130_fd_sc_hd__nor2_2 _35895_ (.A(_07914_),
    .B(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__and2_2 _35896_ (.A(_07914_),
    .B(_07915_),
    .X(_07917_));
 sky130_fd_sc_hd__nor2_2 _35897_ (.A(_07916_),
    .B(_07917_),
    .Y(_07918_));
 sky130_fd_sc_hd__or4_4 _35898_ (.A(_06925_),
    .B(_07434_),
    .C(_07684_),
    .D(_07685_),
    .X(_07919_));
 sky130_fd_sc_hd__and3_2 _35899_ (.A(_06363_),
    .B(_06364_),
    .C(_06653_),
    .X(_07920_));
 sky130_fd_sc_hd__or4b_4 _35900_ (.A(_05767_),
    .B(_07202_),
    .C(_07919_),
    .D_N(_07920_),
    .X(_07921_));
 sky130_fd_sc_hd__nand3_2 _35901_ (.A(_06363_),
    .B(_06368_),
    .C(_06653_),
    .Y(_07922_));
 sky130_fd_sc_hd__a211o_2 _35902_ (.A1(_06929_),
    .A2(_07922_),
    .B1(_07919_),
    .C1(_07202_),
    .X(_07923_));
 sky130_fd_sc_hd__or3_2 _35903_ (.A(_07434_),
    .B(_07684_),
    .C(_07685_),
    .X(_07925_));
 sky130_fd_sc_hd__o21ba_2 _35904_ (.A1(_07445_),
    .A2(_07684_),
    .B1_N(_07685_),
    .X(_07926_));
 sky130_fd_sc_hd__o21a_2 _35905_ (.A1(_07436_),
    .A2(_07925_),
    .B1(_07926_),
    .X(_07927_));
 sky130_fd_sc_hd__and3_2 _35906_ (.A(_07921_),
    .B(_07923_),
    .C(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__xnor2_2 _35907_ (.A(_07918_),
    .B(_07928_),
    .Y(_07929_));
 sky130_fd_sc_hd__nand2_2 _35908_ (.A(_15807_),
    .B(_07929_),
    .Y(_07930_));
 sky130_fd_sc_hd__or2_2 _35909_ (.A(_15807_),
    .B(_07929_),
    .X(_07931_));
 sky130_fd_sc_hd__and2_2 _35910_ (.A(_07930_),
    .B(_07931_),
    .X(_07932_));
 sky130_fd_sc_hd__nor2_2 _35911_ (.A(_07441_),
    .B(_07688_),
    .Y(_07933_));
 sky130_fd_sc_hd__and2_2 _35912_ (.A(_06372_),
    .B(_06658_),
    .X(_07934_));
 sky130_fd_sc_hd__and3_2 _35913_ (.A(_05771_),
    .B(_06075_),
    .C(_07934_),
    .X(_07936_));
 sky130_fd_sc_hd__and4_2 _35914_ (.A(_06936_),
    .B(_07207_),
    .C(_07933_),
    .D(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__a21o_2 _35915_ (.A1(_06078_),
    .A2(_07934_),
    .B1(_06937_),
    .X(_07938_));
 sky130_fd_sc_hd__and3_2 _35916_ (.A(_06936_),
    .B(_07207_),
    .C(_07933_),
    .X(_07939_));
 sky130_fd_sc_hd__or2b_2 _35917_ (.A(_07687_),
    .B_N(_15351_),
    .X(_07940_));
 sky130_fd_sc_hd__nand2_2 _35918_ (.A(_07439_),
    .B(_07940_),
    .Y(_07941_));
 sky130_fd_sc_hd__or2b_2 _35919_ (.A(_15351_),
    .B_N(_07687_),
    .X(_07942_));
 sky130_fd_sc_hd__a22o_2 _35920_ (.A1(_07443_),
    .A2(_07933_),
    .B1(_07941_),
    .B2(_07942_),
    .X(_07943_));
 sky130_fd_sc_hd__a221o_2 _35921_ (.A1(_05781_),
    .A2(_07937_),
    .B1(_07938_),
    .B2(_07939_),
    .C1(_07943_),
    .X(_07944_));
 sky130_fd_sc_hd__a31oi_2 _35922_ (.A1(_03689_),
    .A2(_05774_),
    .A3(_07937_),
    .B1(_07944_),
    .Y(_07945_));
 sky130_fd_sc_hd__xnor2_2 _35923_ (.A(_07932_),
    .B(_07945_),
    .Y(oO[80]));
 sky130_fd_sc_hd__and2b_2 _35924_ (.A_N(_07945_),
    .B(_07932_),
    .X(_07947_));
 sky130_fd_sc_hd__a21oi_2 _35925_ (.A1(_15807_),
    .A2(_07929_),
    .B1(_07947_),
    .Y(_07948_));
 sky130_fd_sc_hd__a21o_2 _35926_ (.A1(_07691_),
    .A2(_07694_),
    .B1(_07807_),
    .X(_07949_));
 sky130_fd_sc_hd__a21oi_2 _35927_ (.A1(_07711_),
    .A2(_07712_),
    .B1(_07709_),
    .Y(_07950_));
 sky130_fd_sc_hd__a2bb2o_2 _35928_ (.A1_N(_16606_),
    .A2_N(_05550_),
    .B1(_03458_),
    .B2(_16614_),
    .X(_07951_));
 sky130_fd_sc_hd__o31a_2 _35929_ (.A1(_04847_),
    .A2(_05550_),
    .A3(_07468_),
    .B1(_07951_),
    .X(_07952_));
 sky130_fd_sc_hd__and2b_2 _35930_ (.A_N(_07950_),
    .B(_07952_),
    .X(_07953_));
 sky130_fd_sc_hd__and2b_2 _35931_ (.A_N(_07952_),
    .B(_07950_),
    .X(_07954_));
 sky130_fd_sc_hd__or2_2 _35932_ (.A(_07953_),
    .B(_07954_),
    .X(_07955_));
 sky130_fd_sc_hd__or4_2 _35933_ (.A(_05980_),
    .B(_05978_),
    .C(_04187_),
    .D(_05231_),
    .X(_07957_));
 sky130_fd_sc_hd__a22o_2 _35934_ (.A1(_06411_),
    .A2(_07472_),
    .B1(_03994_),
    .B2(_06414_),
    .X(_07958_));
 sky130_fd_sc_hd__nand2_2 _35935_ (.A(_07957_),
    .B(_07958_),
    .Y(_07959_));
 sky130_fd_sc_hd__nand2_2 _35936_ (.A(_03345_),
    .B(_07461_),
    .Y(_07960_));
 sky130_fd_sc_hd__xnor2_2 _35937_ (.A(_07959_),
    .B(_07960_),
    .Y(_07961_));
 sky130_fd_sc_hd__nor2_2 _35938_ (.A(_07955_),
    .B(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__and2_2 _35939_ (.A(_07955_),
    .B(_07961_),
    .X(_07963_));
 sky130_fd_sc_hd__nor2_2 _35940_ (.A(_07962_),
    .B(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__and3_2 _35941_ (.A(_07217_),
    .B(_07721_),
    .C(_07964_),
    .X(_07965_));
 sky130_fd_sc_hd__a21oi_2 _35942_ (.A1(_07217_),
    .A2(_07721_),
    .B1(_07964_),
    .Y(_07966_));
 sky130_fd_sc_hd__or2_2 _35943_ (.A(_07965_),
    .B(_07966_),
    .X(_07968_));
 sky130_fd_sc_hd__o22a_2 _35944_ (.A1(_03389_),
    .A2(_04181_),
    .B1(_04901_),
    .B2(_01804_),
    .X(_07969_));
 sky130_fd_sc_hd__a21o_2 _35945_ (.A1(_05533_),
    .A2(_03373_),
    .B1(_07969_),
    .X(_07970_));
 sky130_fd_sc_hd__o21a_2 _35946_ (.A1(_02468_),
    .A2(_06399_),
    .B1(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__a311oi_2 _35947_ (.A1(_06785_),
    .A2(_06789_),
    .A3(_06949_),
    .B1(_07214_),
    .C1(_06947_),
    .Y(_07972_));
 sky130_fd_sc_hd__nand2_2 _35948_ (.A(_07212_),
    .B(_07491_),
    .Y(_07973_));
 sky130_fd_sc_hd__nor2_2 _35949_ (.A(_07698_),
    .B(_07970_),
    .Y(_07974_));
 sky130_fd_sc_hd__o211a_2 _35950_ (.A1(_07972_),
    .A2(_07973_),
    .B1(_07974_),
    .C1(_07493_),
    .X(_07975_));
 sky130_fd_sc_hd__nor3_2 _35951_ (.A(_02468_),
    .B(_06399_),
    .C(_07970_),
    .Y(_07976_));
 sky130_fd_sc_hd__a211o_2 _35952_ (.A1(_07699_),
    .A2(_07971_),
    .B1(_07975_),
    .C1(_07976_),
    .X(_07977_));
 sky130_fd_sc_hd__xor2_2 _35953_ (.A(_07968_),
    .B(_07977_),
    .X(_07979_));
 sky130_fd_sc_hd__xnor2_2 _35954_ (.A(_07730_),
    .B(_07979_),
    .Y(_07980_));
 sky130_fd_sc_hd__a32o_2 _35955_ (.A1(_07769_),
    .A2(_07771_),
    .A3(_07775_),
    .B1(_07776_),
    .B2(_07753_),
    .X(_07981_));
 sky130_fd_sc_hd__and2b_2 _35956_ (.A_N(_07722_),
    .B(_07724_),
    .X(_07982_));
 sky130_fd_sc_hd__buf_1 _35957_ (.A(_05441_),
    .X(_07983_));
 sky130_fd_sc_hd__o31a_2 _35958_ (.A1(_03389_),
    .A2(_07983_),
    .A3(_07736_),
    .B1(_07734_),
    .X(_07984_));
 sky130_fd_sc_hd__nand2_2 _35959_ (.A(_03024_),
    .B(_02928_),
    .Y(_07985_));
 sky130_fd_sc_hd__or3_2 _35960_ (.A(_05983_),
    .B(_07252_),
    .C(_07985_),
    .X(_07986_));
 sky130_fd_sc_hd__o21ai_2 _35961_ (.A1(_05983_),
    .A2(_07252_),
    .B1(_07985_),
    .Y(_07987_));
 sky130_fd_sc_hd__nand2_2 _35962_ (.A(_07986_),
    .B(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__nor2_2 _35963_ (.A(_04504_),
    .B(_05440_),
    .Y(_07990_));
 sky130_fd_sc_hd__xnor2_2 _35964_ (.A(_07988_),
    .B(_07990_),
    .Y(_07991_));
 sky130_fd_sc_hd__nand2_2 _35965_ (.A(_00662_),
    .B(_01757_),
    .Y(_07992_));
 sky130_fd_sc_hd__xnor2_2 _35966_ (.A(_07740_),
    .B(_07992_),
    .Y(_07993_));
 sky130_fd_sc_hd__or3_2 _35967_ (.A(_05979_),
    .B(_00943_),
    .C(_07993_),
    .X(_07994_));
 sky130_fd_sc_hd__o21ai_2 _35968_ (.A1(_05979_),
    .A2(_00944_),
    .B1(_07993_),
    .Y(_07995_));
 sky130_fd_sc_hd__nand2_2 _35969_ (.A(_07994_),
    .B(_07995_),
    .Y(_07996_));
 sky130_fd_sc_hd__o22a_2 _35970_ (.A1(_07511_),
    .A2(_07740_),
    .B1(_07741_),
    .B2(_07743_),
    .X(_07997_));
 sky130_fd_sc_hd__nor2_2 _35971_ (.A(_07996_),
    .B(_07997_),
    .Y(_07998_));
 sky130_fd_sc_hd__and2_2 _35972_ (.A(_07996_),
    .B(_07997_),
    .X(_07999_));
 sky130_fd_sc_hd__nor2_2 _35973_ (.A(_07998_),
    .B(_07999_),
    .Y(_08001_));
 sky130_fd_sc_hd__xnor2_2 _35974_ (.A(_07991_),
    .B(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__a21o_2 _35975_ (.A1(_07739_),
    .A2(_07749_),
    .B1(_07746_),
    .X(_08003_));
 sky130_fd_sc_hd__xnor2_2 _35976_ (.A(_08002_),
    .B(_08003_),
    .Y(_08004_));
 sky130_fd_sc_hd__xnor2_2 _35977_ (.A(_07984_),
    .B(_08004_),
    .Y(_08005_));
 sky130_fd_sc_hd__or2b_2 _35978_ (.A(_07764_),
    .B_N(_07758_),
    .X(_08006_));
 sky130_fd_sc_hd__nand2_2 _35979_ (.A(_07757_),
    .B(_07765_),
    .Y(_08007_));
 sky130_fd_sc_hd__o21ai_2 _35980_ (.A1(_07762_),
    .A2(_07763_),
    .B1(_07760_),
    .Y(_08008_));
 sky130_fd_sc_hd__nand2_2 _35981_ (.A(_07702_),
    .B(_07706_),
    .Y(_08009_));
 sky130_fd_sc_hd__and4_2 _35982_ (.A(_18328_),
    .B(_06488_),
    .C(_01862_),
    .D(_02629_),
    .X(_08010_));
 sky130_fd_sc_hd__o22a_2 _35983_ (.A1(_18344_),
    .A2(_04162_),
    .B1(_05227_),
    .B2(_06491_),
    .X(_08012_));
 sky130_fd_sc_hd__or2_2 _35984_ (.A(_08010_),
    .B(_08012_),
    .X(_08013_));
 sky130_fd_sc_hd__nand2_2 _35985_ (.A(_04138_),
    .B(_04469_),
    .Y(_08014_));
 sky130_fd_sc_hd__xnor2_2 _35986_ (.A(_08013_),
    .B(_08014_),
    .Y(_08015_));
 sky130_fd_sc_hd__xor2_2 _35987_ (.A(_08009_),
    .B(_08015_),
    .X(_08016_));
 sky130_fd_sc_hd__xor2_2 _35988_ (.A(_08008_),
    .B(_08016_),
    .X(_08017_));
 sky130_fd_sc_hd__a21oi_2 _35989_ (.A1(_07716_),
    .A2(_07719_),
    .B1(_08017_),
    .Y(_08018_));
 sky130_fd_sc_hd__and3_2 _35990_ (.A(_07716_),
    .B(_07719_),
    .C(_08017_),
    .X(_08019_));
 sky130_fd_sc_hd__a211o_2 _35991_ (.A1(_08006_),
    .A2(_08007_),
    .B1(_08018_),
    .C1(_08019_),
    .X(_08020_));
 sky130_fd_sc_hd__inv_2 _35992_ (.A(_08020_),
    .Y(_08021_));
 sky130_fd_sc_hd__o211a_2 _35993_ (.A1(_08018_),
    .A2(_08019_),
    .B1(_08006_),
    .C1(_08007_),
    .X(_08023_));
 sky130_fd_sc_hd__a211o_2 _35994_ (.A1(_07767_),
    .A2(_07769_),
    .B1(_08021_),
    .C1(_08023_),
    .X(_08024_));
 sky130_fd_sc_hd__o211ai_2 _35995_ (.A1(_08021_),
    .A2(_08023_),
    .B1(_07767_),
    .C1(_07769_),
    .Y(_08025_));
 sky130_fd_sc_hd__nand3_2 _35996_ (.A(_08005_),
    .B(_08024_),
    .C(_08025_),
    .Y(_08026_));
 sky130_fd_sc_hd__a21o_2 _35997_ (.A1(_08024_),
    .A2(_08025_),
    .B1(_08005_),
    .X(_08027_));
 sky130_fd_sc_hd__and3_2 _35998_ (.A(_07982_),
    .B(_08026_),
    .C(_08027_),
    .X(_08028_));
 sky130_fd_sc_hd__a21oi_2 _35999_ (.A1(_08026_),
    .A2(_08027_),
    .B1(_07982_),
    .Y(_08029_));
 sky130_fd_sc_hd__nor2_2 _36000_ (.A(_08028_),
    .B(_08029_),
    .Y(_08030_));
 sky130_fd_sc_hd__xor2_2 _36001_ (.A(_07981_),
    .B(_08030_),
    .X(_08031_));
 sky130_fd_sc_hd__xnor2_2 _36002_ (.A(_07980_),
    .B(_08031_),
    .Y(_08032_));
 sky130_fd_sc_hd__and2_2 _36003_ (.A(_07729_),
    .B(_07780_),
    .X(_08034_));
 sky130_fd_sc_hd__xnor2_2 _36004_ (.A(_08032_),
    .B(_08034_),
    .Y(_08035_));
 sky130_fd_sc_hd__nand2_2 _36005_ (.A(_07732_),
    .B(_07778_),
    .Y(_08036_));
 sky130_fd_sc_hd__o31a_2 _36006_ (.A1(_07484_),
    .A2(_07486_),
    .A3(_07777_),
    .B1(_08036_),
    .X(_08037_));
 sky130_fd_sc_hd__and2b_2 _36007_ (.A_N(_07750_),
    .B(_07751_),
    .X(_08038_));
 sky130_fd_sc_hd__and2b_2 _36008_ (.A_N(_07733_),
    .B(_07752_),
    .X(_08039_));
 sky130_fd_sc_hd__nor2_2 _36009_ (.A(_08038_),
    .B(_08039_),
    .Y(_08040_));
 sky130_fd_sc_hd__xnor2_2 _36010_ (.A(_08037_),
    .B(_08040_),
    .Y(_08041_));
 sky130_fd_sc_hd__nor2_2 _36011_ (.A(_08035_),
    .B(_08041_),
    .Y(_08042_));
 sky130_fd_sc_hd__and2_2 _36012_ (.A(_08035_),
    .B(_08041_),
    .X(_08043_));
 sky130_fd_sc_hd__nor2_2 _36013_ (.A(_08042_),
    .B(_08043_),
    .Y(_08045_));
 sky130_fd_sc_hd__nor2_2 _36014_ (.A(_07783_),
    .B(_07794_),
    .Y(_08046_));
 sky130_fd_sc_hd__xnor2_2 _36015_ (.A(_08045_),
    .B(_08046_),
    .Y(_08047_));
 sky130_fd_sc_hd__xnor2_2 _36016_ (.A(_07790_),
    .B(_08047_),
    .Y(_08048_));
 sky130_fd_sc_hd__nand2_2 _36017_ (.A(_07796_),
    .B(_07799_),
    .Y(_08049_));
 sky130_fd_sc_hd__xor2_2 _36018_ (.A(_08048_),
    .B(_08049_),
    .X(_08050_));
 sky130_fd_sc_hd__a21o_2 _36019_ (.A1(_07805_),
    .A2(_07949_),
    .B1(_08050_),
    .X(_08051_));
 sky130_fd_sc_hd__nand3_2 _36020_ (.A(_07805_),
    .B(_07949_),
    .C(_08050_),
    .Y(_08052_));
 sky130_fd_sc_hd__nand2_2 _36021_ (.A(_08051_),
    .B(_08052_),
    .Y(_08053_));
 sky130_fd_sc_hd__and2_2 _36022_ (.A(_07895_),
    .B(_07896_),
    .X(_08054_));
 sky130_fd_sc_hd__and4_2 _36023_ (.A(iY[53]),
    .B(iY[54]),
    .C(iX[59]),
    .D(iX[60]),
    .X(_08056_));
 sky130_fd_sc_hd__a22oi_2 _36024_ (.A1(iY[54]),
    .A2(iX[59]),
    .B1(iX[60]),
    .B2(iY[53]),
    .Y(_08057_));
 sky130_fd_sc_hd__nand2_2 _36025_ (.A(iY[55]),
    .B(iX[58]),
    .Y(_08058_));
 sky130_fd_sc_hd__o21a_2 _36026_ (.A1(_08056_),
    .A2(_08057_),
    .B1(_08058_),
    .X(_08059_));
 sky130_fd_sc_hd__nor3_2 _36027_ (.A(_08056_),
    .B(_08057_),
    .C(_08058_),
    .Y(_08060_));
 sky130_fd_sc_hd__nor2_2 _36028_ (.A(_08059_),
    .B(_08060_),
    .Y(_08061_));
 sky130_fd_sc_hd__inv_2 _36029_ (.A(_08061_),
    .Y(_08062_));
 sky130_fd_sc_hd__nand2_2 _36030_ (.A(iY[50]),
    .B(iX[63]),
    .Y(_08063_));
 sky130_fd_sc_hd__xnor2_2 _36031_ (.A(_07820_),
    .B(_08063_),
    .Y(_08064_));
 sky130_fd_sc_hd__and2_2 _36032_ (.A(iY[52]),
    .B(iX[61]),
    .X(_08065_));
 sky130_fd_sc_hd__nor2_2 _36033_ (.A(_08064_),
    .B(_08065_),
    .Y(_08067_));
 sky130_fd_sc_hd__and2_2 _36034_ (.A(_08064_),
    .B(_08065_),
    .X(_08068_));
 sky130_fd_sc_hd__nor2_2 _36035_ (.A(_08067_),
    .B(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__o21a_2 _36036_ (.A1(_07821_),
    .A2(_07826_),
    .B1(_08069_),
    .X(_08070_));
 sky130_fd_sc_hd__nor3_2 _36037_ (.A(_07821_),
    .B(_07826_),
    .C(_08069_),
    .Y(_08071_));
 sky130_fd_sc_hd__or2_2 _36038_ (.A(_08070_),
    .B(_08071_),
    .X(_08072_));
 sky130_fd_sc_hd__nor2_2 _36039_ (.A(_08062_),
    .B(_08072_),
    .Y(_08073_));
 sky130_fd_sc_hd__and2_2 _36040_ (.A(_08062_),
    .B(_08072_),
    .X(_08074_));
 sky130_fd_sc_hd__or2_2 _36041_ (.A(_08073_),
    .B(_08074_),
    .X(_08075_));
 sky130_fd_sc_hd__or3_2 _36042_ (.A(_07580_),
    .B(_07581_),
    .C(_08075_),
    .X(_08076_));
 sky130_fd_sc_hd__o21ai_2 _36043_ (.A1(_07580_),
    .A2(_07581_),
    .B1(_08075_),
    .Y(_08077_));
 sky130_fd_sc_hd__nand2_2 _36044_ (.A(_08076_),
    .B(_08077_),
    .Y(_08078_));
 sky130_fd_sc_hd__a31o_2 _36045_ (.A1(_07583_),
    .A2(_07585_),
    .A3(_07812_),
    .B1(_07833_),
    .X(_08079_));
 sky130_fd_sc_hd__and2b_2 _36046_ (.A_N(_08078_),
    .B(_08079_),
    .X(_08080_));
 sky130_fd_sc_hd__and2b_2 _36047_ (.A_N(_08079_),
    .B(_08078_),
    .X(_08081_));
 sky130_fd_sc_hd__or2_2 _36048_ (.A(_08080_),
    .B(_08081_),
    .X(_08082_));
 sky130_fd_sc_hd__or2b_2 _36049_ (.A(_07844_),
    .B_N(_07843_),
    .X(_08083_));
 sky130_fd_sc_hd__and4_2 _36050_ (.A(iX[53]),
    .B(iX[54]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_08084_));
 sky130_fd_sc_hd__a22oi_2 _36051_ (.A1(iX[54]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[53]),
    .Y(_08085_));
 sky130_fd_sc_hd__nor2_2 _36052_ (.A(_08084_),
    .B(_08085_),
    .Y(_08086_));
 sky130_fd_sc_hd__nand2_2 _36053_ (.A(iX[52]),
    .B(iY[61]),
    .Y(_08088_));
 sky130_fd_sc_hd__xnor2_2 _36054_ (.A(_08086_),
    .B(_08088_),
    .Y(_08089_));
 sky130_fd_sc_hd__o21ba_2 _36055_ (.A1(_07840_),
    .A2(_07842_),
    .B1_N(_07839_),
    .X(_08090_));
 sky130_fd_sc_hd__xnor2_2 _36056_ (.A(_08089_),
    .B(_08090_),
    .Y(_08091_));
 sky130_fd_sc_hd__nand2_2 _36057_ (.A(iX[51]),
    .B(iY[62]),
    .Y(_08092_));
 sky130_fd_sc_hd__xor2_2 _36058_ (.A(_08091_),
    .B(_08092_),
    .X(_08093_));
 sky130_fd_sc_hd__a21oi_2 _36059_ (.A1(_08083_),
    .A2(_07849_),
    .B1(_08093_),
    .Y(_08094_));
 sky130_fd_sc_hd__and3_2 _36060_ (.A(_08083_),
    .B(_07849_),
    .C(_08093_),
    .X(_08095_));
 sky130_fd_sc_hd__nor2_2 _36061_ (.A(_08094_),
    .B(_08095_),
    .Y(_08096_));
 sky130_fd_sc_hd__a21oi_2 _36062_ (.A1(iX[50]),
    .A2(iY[63]),
    .B1(_08096_),
    .Y(_08097_));
 sky130_fd_sc_hd__and3_2 _36063_ (.A(iX[50]),
    .B(iY[63]),
    .C(_08096_),
    .X(_08099_));
 sky130_fd_sc_hd__nor2_2 _36064_ (.A(_08097_),
    .B(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__or2b_2 _36065_ (.A(_07864_),
    .B_N(_07870_),
    .X(_08101_));
 sky130_fd_sc_hd__or2b_2 _36066_ (.A(_07863_),
    .B_N(_07871_),
    .X(_08102_));
 sky130_fd_sc_hd__and2b_2 _36067_ (.A_N(_07828_),
    .B(_07827_),
    .X(_08103_));
 sky130_fd_sc_hd__o21ba_2 _36068_ (.A1(_07866_),
    .A2(_07868_),
    .B1_N(_07865_),
    .X(_08104_));
 sky130_fd_sc_hd__o21ba_2 _36069_ (.A1(_07816_),
    .A2(_07818_),
    .B1_N(_07815_),
    .X(_08105_));
 sky130_fd_sc_hd__and4_2 _36070_ (.A(iX[56]),
    .B(iY[56]),
    .C(iX[57]),
    .D(iY[57]),
    .X(_08106_));
 sky130_fd_sc_hd__a22oi_2 _36071_ (.A1(iY[56]),
    .A2(iX[57]),
    .B1(iY[57]),
    .B2(iX[56]),
    .Y(_08107_));
 sky130_fd_sc_hd__nor2_2 _36072_ (.A(_08106_),
    .B(_08107_),
    .Y(_08108_));
 sky130_fd_sc_hd__nand2_2 _36073_ (.A(iX[55]),
    .B(iY[58]),
    .Y(_08110_));
 sky130_fd_sc_hd__xnor2_2 _36074_ (.A(_08108_),
    .B(_08110_),
    .Y(_08111_));
 sky130_fd_sc_hd__xnor2_2 _36075_ (.A(_08105_),
    .B(_08111_),
    .Y(_08112_));
 sky130_fd_sc_hd__xnor2_2 _36076_ (.A(_08104_),
    .B(_08112_),
    .Y(_08113_));
 sky130_fd_sc_hd__o21a_2 _36077_ (.A1(_08103_),
    .A2(_07830_),
    .B1(_08113_),
    .X(_08114_));
 sky130_fd_sc_hd__nor3_2 _36078_ (.A(_08103_),
    .B(_07830_),
    .C(_08113_),
    .Y(_08115_));
 sky130_fd_sc_hd__a211oi_2 _36079_ (.A1(_08101_),
    .A2(_08102_),
    .B1(_08114_),
    .C1(_08115_),
    .Y(_08116_));
 sky130_fd_sc_hd__o211a_2 _36080_ (.A1(_08114_),
    .A2(_08115_),
    .B1(_08101_),
    .C1(_08102_),
    .X(_08117_));
 sky130_fd_sc_hd__nor2_2 _36081_ (.A(_07873_),
    .B(_07875_),
    .Y(_08118_));
 sky130_fd_sc_hd__or3_2 _36082_ (.A(_08116_),
    .B(_08117_),
    .C(_08118_),
    .X(_08119_));
 sky130_fd_sc_hd__o21ai_2 _36083_ (.A1(_08116_),
    .A2(_08117_),
    .B1(_08118_),
    .Y(_08121_));
 sky130_fd_sc_hd__and3_2 _36084_ (.A(_08100_),
    .B(_08119_),
    .C(_08121_),
    .X(_08122_));
 sky130_fd_sc_hd__a21oi_2 _36085_ (.A1(_08119_),
    .A2(_08121_),
    .B1(_08100_),
    .Y(_08123_));
 sky130_fd_sc_hd__nor3_2 _36086_ (.A(_07835_),
    .B(_08122_),
    .C(_08123_),
    .Y(_08124_));
 sky130_fd_sc_hd__o21a_2 _36087_ (.A1(_08122_),
    .A2(_08123_),
    .B1(_07835_),
    .X(_08125_));
 sky130_fd_sc_hd__or2_2 _36088_ (.A(_08124_),
    .B(_08125_),
    .X(_08126_));
 sky130_fd_sc_hd__a21oi_2 _36089_ (.A1(_07878_),
    .A2(_07881_),
    .B1(_08126_),
    .Y(_08127_));
 sky130_fd_sc_hd__and3_2 _36090_ (.A(_07878_),
    .B(_07881_),
    .C(_08126_),
    .X(_08128_));
 sky130_fd_sc_hd__or3_2 _36091_ (.A(_08082_),
    .B(_08127_),
    .C(_08128_),
    .X(_08129_));
 sky130_fd_sc_hd__o21ai_2 _36092_ (.A1(_08127_),
    .A2(_08128_),
    .B1(_08082_),
    .Y(_08130_));
 sky130_fd_sc_hd__and3_2 _36093_ (.A(_07888_),
    .B(_08129_),
    .C(_08130_),
    .X(_08132_));
 sky130_fd_sc_hd__a21oi_2 _36094_ (.A1(_08129_),
    .A2(_08130_),
    .B1(_07888_),
    .Y(_08133_));
 sky130_fd_sc_hd__a211oi_2 _36095_ (.A1(_07883_),
    .A2(_07886_),
    .B1(_08132_),
    .C1(_08133_),
    .Y(_08134_));
 sky130_fd_sc_hd__o211a_2 _36096_ (.A1(_08132_),
    .A2(_08133_),
    .B1(_07883_),
    .C1(_07886_),
    .X(_08135_));
 sky130_fd_sc_hd__a211oi_2 _36097_ (.A1(_07890_),
    .A2(_07893_),
    .B1(_08134_),
    .C1(_08135_),
    .Y(_08136_));
 sky130_fd_sc_hd__o211a_2 _36098_ (.A1(_08134_),
    .A2(_08135_),
    .B1(_07890_),
    .C1(_07893_),
    .X(_08137_));
 sky130_fd_sc_hd__a211oi_2 _36099_ (.A1(_07852_),
    .A2(_07857_),
    .B1(_08136_),
    .C1(_08137_),
    .Y(_08138_));
 sky130_fd_sc_hd__o211a_2 _36100_ (.A1(_08136_),
    .A2(_08137_),
    .B1(_07852_),
    .C1(_07857_),
    .X(_08139_));
 sky130_fd_sc_hd__nor2_2 _36101_ (.A(_08138_),
    .B(_08139_),
    .Y(_08140_));
 sky130_fd_sc_hd__o21a_2 _36102_ (.A1(_08054_),
    .A2(_07898_),
    .B1(_08140_),
    .X(_08141_));
 sky130_fd_sc_hd__nor3_2 _36103_ (.A(_08054_),
    .B(_07898_),
    .C(_08140_),
    .Y(_08143_));
 sky130_fd_sc_hd__or2_2 _36104_ (.A(_08141_),
    .B(_08143_),
    .X(_08144_));
 sky130_fd_sc_hd__o21bai_2 _36105_ (.A1(_07905_),
    .A2(_07910_),
    .B1_N(_07903_),
    .Y(_08145_));
 sky130_fd_sc_hd__xnor2_2 _36106_ (.A(_08144_),
    .B(_08145_),
    .Y(_08146_));
 sky130_fd_sc_hd__xor2_2 _36107_ (.A(_08053_),
    .B(_08146_),
    .X(_08147_));
 sky130_fd_sc_hd__xnor2_2 _36108_ (.A(_16134_),
    .B(_08147_),
    .Y(_08148_));
 sky130_fd_sc_hd__or2b_2 _36109_ (.A(_15575_),
    .B_N(_07912_),
    .X(_08149_));
 sky130_fd_sc_hd__o31a_2 _36110_ (.A1(_07808_),
    .A2(_07809_),
    .A3(_07911_),
    .B1(_08149_),
    .X(_08150_));
 sky130_fd_sc_hd__xor2_2 _36111_ (.A(_08148_),
    .B(_08150_),
    .X(_08151_));
 sky130_fd_sc_hd__and2b_2 _36112_ (.A_N(_07928_),
    .B(_07918_),
    .X(_08152_));
 sky130_fd_sc_hd__nor2_2 _36113_ (.A(_07916_),
    .B(_08152_),
    .Y(_08154_));
 sky130_fd_sc_hd__xnor2_2 _36114_ (.A(_08151_),
    .B(_08154_),
    .Y(_08155_));
 sky130_fd_sc_hd__and2b_2 _36115_ (.A_N(_08155_),
    .B(_16034_),
    .X(_08156_));
 sky130_fd_sc_hd__or2b_2 _36116_ (.A(_16034_),
    .B_N(_08155_),
    .X(_08157_));
 sky130_fd_sc_hd__and2b_2 _36117_ (.A_N(_08156_),
    .B(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__xnor2_2 _36118_ (.A(_07948_),
    .B(_08158_),
    .Y(oO[81]));
 sky130_fd_sc_hd__or2b_2 _36119_ (.A(_08048_),
    .B_N(_08049_),
    .X(_08159_));
 sky130_fd_sc_hd__nor2_2 _36120_ (.A(_08037_),
    .B(_08040_),
    .Y(_08160_));
 sky130_fd_sc_hd__or2_2 _36121_ (.A(_07968_),
    .B(_07977_),
    .X(_08161_));
 sky130_fd_sc_hd__a21o_2 _36122_ (.A1(_05533_),
    .A2(_03373_),
    .B1(_07976_),
    .X(_08162_));
 sky130_fd_sc_hd__buf_1 _36123_ (.A(_04901_),
    .X(_08164_));
 sky130_fd_sc_hd__o22a_2 _36124_ (.A1(_04504_),
    .A2(_06786_),
    .B1(_08164_),
    .B2(_16606_),
    .X(_08165_));
 sky130_fd_sc_hd__a21oi_2 _36125_ (.A1(_05533_),
    .A2(_03938_),
    .B1(_08165_),
    .Y(_08166_));
 sky130_fd_sc_hd__o21ai_2 _36126_ (.A1(_07975_),
    .A2(_08162_),
    .B1(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__or3_2 _36127_ (.A(_07975_),
    .B(_08166_),
    .C(_08162_),
    .X(_08168_));
 sky130_fd_sc_hd__and2_2 _36128_ (.A(_08167_),
    .B(_08168_),
    .X(_08169_));
 sky130_fd_sc_hd__or4_2 _36129_ (.A(_05980_),
    .B(_05978_),
    .C(_05231_),
    .D(_06797_),
    .X(_08170_));
 sky130_fd_sc_hd__a22o_2 _36130_ (.A1(_06411_),
    .A2(_03994_),
    .B1(_03458_),
    .B2(_06414_),
    .X(_08171_));
 sky130_fd_sc_hd__and2_2 _36131_ (.A(_08170_),
    .B(_08171_),
    .X(_08172_));
 sky130_fd_sc_hd__nor2_2 _36132_ (.A(_05500_),
    .B(_06023_),
    .Y(_08173_));
 sky130_fd_sc_hd__xnor2_2 _36133_ (.A(_08172_),
    .B(_08173_),
    .Y(_08175_));
 sky130_fd_sc_hd__and3_2 _36134_ (.A(_16614_),
    .B(_06783_),
    .C(_07468_),
    .X(_08176_));
 sky130_fd_sc_hd__xnor2_2 _36135_ (.A(_08175_),
    .B(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__xnor2_2 _36136_ (.A(_08169_),
    .B(_08177_),
    .Y(_08178_));
 sky130_fd_sc_hd__xnor2_2 _36137_ (.A(_08161_),
    .B(_08178_),
    .Y(_08179_));
 sky130_fd_sc_hd__o31a_2 _36138_ (.A1(_04504_),
    .A2(_05441_),
    .A3(_07988_),
    .B1(_07986_),
    .X(_08180_));
 sky130_fd_sc_hd__nor2_2 _36139_ (.A(_04501_),
    .B(_05931_),
    .Y(_08181_));
 sky130_fd_sc_hd__and3_2 _36140_ (.A(_05507_),
    .B(_02928_),
    .C(_08181_),
    .X(_08182_));
 sky130_fd_sc_hd__a21oi_2 _36141_ (.A1(_05507_),
    .A2(_04781_),
    .B1(_08181_),
    .Y(_08183_));
 sky130_fd_sc_hd__nor2_2 _36142_ (.A(_08182_),
    .B(_08183_),
    .Y(_08184_));
 sky130_fd_sc_hd__nor2_2 _36143_ (.A(_05983_),
    .B(_05440_),
    .Y(_08186_));
 sky130_fd_sc_hd__xor2_2 _36144_ (.A(_08184_),
    .B(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__nand2_2 _36145_ (.A(_04138_),
    .B(_00567_),
    .Y(_08188_));
 sky130_fd_sc_hd__o22a_2 _36146_ (.A1(_05522_),
    .A2(_07259_),
    .B1(_02311_),
    .B2(_05504_),
    .X(_08189_));
 sky130_fd_sc_hd__o21bai_2 _36147_ (.A1(_07992_),
    .A2(_08188_),
    .B1_N(_08189_),
    .Y(_08190_));
 sky130_fd_sc_hd__nand2_2 _36148_ (.A(_03973_),
    .B(_03327_),
    .Y(_08191_));
 sky130_fd_sc_hd__xnor2_2 _36149_ (.A(_08190_),
    .B(_08191_),
    .Y(_08192_));
 sky130_fd_sc_hd__o21a_2 _36150_ (.A1(_07740_),
    .A2(_07992_),
    .B1(_07994_),
    .X(_08193_));
 sky130_fd_sc_hd__or2_2 _36151_ (.A(_08192_),
    .B(_08193_),
    .X(_08194_));
 sky130_fd_sc_hd__nand2_2 _36152_ (.A(_08192_),
    .B(_08193_),
    .Y(_08195_));
 sky130_fd_sc_hd__and2_2 _36153_ (.A(_08194_),
    .B(_08195_),
    .X(_08197_));
 sky130_fd_sc_hd__nand2_2 _36154_ (.A(_08187_),
    .B(_08197_),
    .Y(_08198_));
 sky130_fd_sc_hd__or2_2 _36155_ (.A(_08187_),
    .B(_08197_),
    .X(_08199_));
 sky130_fd_sc_hd__nand2_2 _36156_ (.A(_08198_),
    .B(_08199_),
    .Y(_08200_));
 sky130_fd_sc_hd__a21o_2 _36157_ (.A1(_07991_),
    .A2(_08001_),
    .B1(_07998_),
    .X(_08201_));
 sky130_fd_sc_hd__xnor2_2 _36158_ (.A(_08200_),
    .B(_08201_),
    .Y(_08202_));
 sky130_fd_sc_hd__xnor2_2 _36159_ (.A(_08180_),
    .B(_08202_),
    .Y(_08203_));
 sky130_fd_sc_hd__a21o_2 _36160_ (.A1(_07716_),
    .A2(_07719_),
    .B1(_08017_),
    .X(_08204_));
 sky130_fd_sc_hd__or2b_2 _36161_ (.A(_08015_),
    .B_N(_08009_),
    .X(_08205_));
 sky130_fd_sc_hd__or2b_2 _36162_ (.A(_08016_),
    .B_N(_08008_),
    .X(_08206_));
 sky130_fd_sc_hd__o21ba_2 _36163_ (.A1(_08012_),
    .A2(_08014_),
    .B1_N(_08010_),
    .X(_08208_));
 sky130_fd_sc_hd__o21ai_2 _36164_ (.A1(_07959_),
    .A2(_07960_),
    .B1(_07957_),
    .Y(_08209_));
 sky130_fd_sc_hd__nand2_2 _36165_ (.A(_18734_),
    .B(_03438_),
    .Y(_08210_));
 sky130_fd_sc_hd__or3_2 _36166_ (.A(_06491_),
    .B(_05227_),
    .C(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__a22o_2 _36167_ (.A1(_06488_),
    .A2(_06983_),
    .B1(_07461_),
    .B2(_18328_),
    .X(_08212_));
 sky130_fd_sc_hd__nand2_2 _36168_ (.A(_08211_),
    .B(_08212_),
    .Y(_08213_));
 sky130_fd_sc_hd__nor2_2 _36169_ (.A(_03341_),
    .B(_06816_),
    .Y(_08214_));
 sky130_fd_sc_hd__xor2_2 _36170_ (.A(_08213_),
    .B(_08214_),
    .X(_08215_));
 sky130_fd_sc_hd__xnor2_2 _36171_ (.A(_08209_),
    .B(_08215_),
    .Y(_08216_));
 sky130_fd_sc_hd__xnor2_2 _36172_ (.A(_08208_),
    .B(_08216_),
    .Y(_08217_));
 sky130_fd_sc_hd__o21ai_2 _36173_ (.A1(_07953_),
    .A2(_07962_),
    .B1(_08217_),
    .Y(_08219_));
 sky130_fd_sc_hd__or3_2 _36174_ (.A(_07953_),
    .B(_07962_),
    .C(_08217_),
    .X(_08220_));
 sky130_fd_sc_hd__nand2_2 _36175_ (.A(_08219_),
    .B(_08220_),
    .Y(_08221_));
 sky130_fd_sc_hd__a21o_2 _36176_ (.A1(_08205_),
    .A2(_08206_),
    .B1(_08221_),
    .X(_08222_));
 sky130_fd_sc_hd__inv_2 _36177_ (.A(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__and3_2 _36178_ (.A(_08205_),
    .B(_08206_),
    .C(_08221_),
    .X(_08224_));
 sky130_fd_sc_hd__a211o_2 _36179_ (.A1(_08204_),
    .A2(_08020_),
    .B1(_08223_),
    .C1(_08224_),
    .X(_08225_));
 sky130_fd_sc_hd__o211ai_2 _36180_ (.A1(_08223_),
    .A2(_08224_),
    .B1(_08204_),
    .C1(_08020_),
    .Y(_08226_));
 sky130_fd_sc_hd__nand3_2 _36181_ (.A(_08203_),
    .B(_08225_),
    .C(_08226_),
    .Y(_08227_));
 sky130_fd_sc_hd__a21o_2 _36182_ (.A1(_08225_),
    .A2(_08226_),
    .B1(_08203_),
    .X(_08228_));
 sky130_fd_sc_hd__and3_2 _36183_ (.A(_07965_),
    .B(_08227_),
    .C(_08228_),
    .X(_08230_));
 sky130_fd_sc_hd__a21oi_2 _36184_ (.A1(_08227_),
    .A2(_08228_),
    .B1(_07965_),
    .Y(_08231_));
 sky130_fd_sc_hd__a211oi_2 _36185_ (.A1(_08024_),
    .A2(_08026_),
    .B1(_08230_),
    .C1(_08231_),
    .Y(_08232_));
 sky130_fd_sc_hd__o211a_2 _36186_ (.A1(_08230_),
    .A2(_08231_),
    .B1(_08024_),
    .C1(_08026_),
    .X(_08233_));
 sky130_fd_sc_hd__or2_2 _36187_ (.A(_08232_),
    .B(_08233_),
    .X(_08234_));
 sky130_fd_sc_hd__xnor2_2 _36188_ (.A(_08179_),
    .B(_08234_),
    .Y(_08235_));
 sky130_fd_sc_hd__nand2_2 _36189_ (.A(_07727_),
    .B(_07979_),
    .Y(_08236_));
 sky130_fd_sc_hd__a21bo_2 _36190_ (.A1(_07980_),
    .A2(_08031_),
    .B1_N(_08236_),
    .X(_08237_));
 sky130_fd_sc_hd__xnor2_2 _36191_ (.A(_08235_),
    .B(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__a21o_2 _36192_ (.A1(_07981_),
    .A2(_08030_),
    .B1(_08028_),
    .X(_08239_));
 sky130_fd_sc_hd__and2b_2 _36193_ (.A_N(_08002_),
    .B(_08003_),
    .X(_08241_));
 sky130_fd_sc_hd__and2b_2 _36194_ (.A_N(_07984_),
    .B(_08004_),
    .X(_08242_));
 sky130_fd_sc_hd__nor2_2 _36195_ (.A(_08241_),
    .B(_08242_),
    .Y(_08243_));
 sky130_fd_sc_hd__xnor2_2 _36196_ (.A(_08239_),
    .B(_08243_),
    .Y(_08244_));
 sky130_fd_sc_hd__xor2_2 _36197_ (.A(_08238_),
    .B(_08244_),
    .X(_08245_));
 sky130_fd_sc_hd__o21ba_2 _36198_ (.A1(_08032_),
    .A2(_08034_),
    .B1_N(_08042_),
    .X(_08246_));
 sky130_fd_sc_hd__xnor2_2 _36199_ (.A(_08245_),
    .B(_08246_),
    .Y(_08247_));
 sky130_fd_sc_hd__xnor2_2 _36200_ (.A(_08160_),
    .B(_08247_),
    .Y(_08248_));
 sky130_fd_sc_hd__and2b_2 _36201_ (.A_N(_08046_),
    .B(_08045_),
    .X(_08249_));
 sky130_fd_sc_hd__a21oi_2 _36202_ (.A1(_07790_),
    .A2(_08047_),
    .B1(_08249_),
    .Y(_08250_));
 sky130_fd_sc_hd__xnor2_2 _36203_ (.A(_08248_),
    .B(_08250_),
    .Y(_08252_));
 sky130_fd_sc_hd__a21o_2 _36204_ (.A1(_08159_),
    .A2(_08051_),
    .B1(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__nand3_2 _36205_ (.A(_08159_),
    .B(_08051_),
    .C(_08252_),
    .Y(_08254_));
 sky130_fd_sc_hd__and3_2 _36206_ (.A(iY[52]),
    .B(iX[63]),
    .C(_07820_),
    .X(_08255_));
 sky130_fd_sc_hd__a22oi_2 _36207_ (.A1(iY[52]),
    .A2(iX[62]),
    .B1(iX[63]),
    .B2(iY[51]),
    .Y(_08256_));
 sky130_fd_sc_hd__or2_2 _36208_ (.A(_08255_),
    .B(_08256_),
    .X(_08257_));
 sky130_fd_sc_hd__a31o_2 _36209_ (.A1(iY[50]),
    .A2(iX[63]),
    .A3(_07820_),
    .B1(_08068_),
    .X(_08258_));
 sky130_fd_sc_hd__xnor2_2 _36210_ (.A(_08257_),
    .B(_08258_),
    .Y(_08259_));
 sky130_fd_sc_hd__and4_2 _36211_ (.A(iY[53]),
    .B(iY[54]),
    .C(iX[60]),
    .D(iX[61]),
    .X(_08260_));
 sky130_fd_sc_hd__a22oi_2 _36212_ (.A1(iY[54]),
    .A2(iX[60]),
    .B1(iX[61]),
    .B2(iY[53]),
    .Y(_08261_));
 sky130_fd_sc_hd__nor2_2 _36213_ (.A(_08260_),
    .B(_08261_),
    .Y(_08263_));
 sky130_fd_sc_hd__nand2_2 _36214_ (.A(iY[55]),
    .B(iX[59]),
    .Y(_08264_));
 sky130_fd_sc_hd__xnor2_2 _36215_ (.A(_08263_),
    .B(_08264_),
    .Y(_08265_));
 sky130_fd_sc_hd__nand2_2 _36216_ (.A(_08259_),
    .B(_08265_),
    .Y(_08266_));
 sky130_fd_sc_hd__or2_2 _36217_ (.A(_08259_),
    .B(_08265_),
    .X(_08267_));
 sky130_fd_sc_hd__nand2_2 _36218_ (.A(_08266_),
    .B(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__or2_2 _36219_ (.A(_08076_),
    .B(_08268_),
    .X(_08269_));
 sky130_fd_sc_hd__nand2_2 _36220_ (.A(_08076_),
    .B(_08268_),
    .Y(_08270_));
 sky130_fd_sc_hd__nand2_2 _36221_ (.A(_08269_),
    .B(_08270_),
    .Y(_08271_));
 sky130_fd_sc_hd__inv_2 _36222_ (.A(_08122_),
    .Y(_08272_));
 sky130_fd_sc_hd__and4_2 _36223_ (.A(iX[54]),
    .B(iX[55]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_08274_));
 sky130_fd_sc_hd__a22oi_2 _36224_ (.A1(iX[55]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[54]),
    .Y(_08275_));
 sky130_fd_sc_hd__nor2_2 _36225_ (.A(_08274_),
    .B(_08275_),
    .Y(_08276_));
 sky130_fd_sc_hd__nand2_2 _36226_ (.A(iX[53]),
    .B(iY[61]),
    .Y(_08277_));
 sky130_fd_sc_hd__xnor2_2 _36227_ (.A(_08276_),
    .B(_08277_),
    .Y(_08278_));
 sky130_fd_sc_hd__o21ba_2 _36228_ (.A1(_08085_),
    .A2(_08088_),
    .B1_N(_08084_),
    .X(_08279_));
 sky130_fd_sc_hd__xnor2_2 _36229_ (.A(_08278_),
    .B(_08279_),
    .Y(_08280_));
 sky130_fd_sc_hd__and2_2 _36230_ (.A(iX[52]),
    .B(iY[62]),
    .X(_08281_));
 sky130_fd_sc_hd__or2_2 _36231_ (.A(_08280_),
    .B(_08281_),
    .X(_08282_));
 sky130_fd_sc_hd__nand2_2 _36232_ (.A(_08280_),
    .B(_08281_),
    .Y(_08283_));
 sky130_fd_sc_hd__and2b_2 _36233_ (.A_N(_08090_),
    .B(_08089_),
    .X(_08285_));
 sky130_fd_sc_hd__a31o_2 _36234_ (.A1(iX[51]),
    .A2(iY[62]),
    .A3(_08091_),
    .B1(_08285_),
    .X(_08286_));
 sky130_fd_sc_hd__nand3_2 _36235_ (.A(_08282_),
    .B(_08283_),
    .C(_08286_),
    .Y(_08287_));
 sky130_fd_sc_hd__a21o_2 _36236_ (.A1(_08282_),
    .A2(_08283_),
    .B1(_08286_),
    .X(_08288_));
 sky130_fd_sc_hd__nand2_2 _36237_ (.A(_08287_),
    .B(_08288_),
    .Y(_08289_));
 sky130_fd_sc_hd__nand2_2 _36238_ (.A(iX[51]),
    .B(iY[63]),
    .Y(_08290_));
 sky130_fd_sc_hd__nand2_2 _36239_ (.A(_08289_),
    .B(_08290_),
    .Y(_08291_));
 sky130_fd_sc_hd__or2_2 _36240_ (.A(_08289_),
    .B(_08290_),
    .X(_08292_));
 sky130_fd_sc_hd__and2_2 _36241_ (.A(_08291_),
    .B(_08292_),
    .X(_08293_));
 sky130_fd_sc_hd__or2b_2 _36242_ (.A(_08105_),
    .B_N(_08111_),
    .X(_08294_));
 sky130_fd_sc_hd__or2b_2 _36243_ (.A(_08104_),
    .B_N(_08112_),
    .X(_08296_));
 sky130_fd_sc_hd__o21ba_2 _36244_ (.A1(_08107_),
    .A2(_08110_),
    .B1_N(_08106_),
    .X(_08297_));
 sky130_fd_sc_hd__and4_2 _36245_ (.A(iY[56]),
    .B(iX[57]),
    .C(iY[57]),
    .D(iX[58]),
    .X(_08298_));
 sky130_fd_sc_hd__a22oi_2 _36246_ (.A1(iX[57]),
    .A2(iY[57]),
    .B1(iX[58]),
    .B2(iY[56]),
    .Y(_08299_));
 sky130_fd_sc_hd__nand2_2 _36247_ (.A(iX[56]),
    .B(iY[58]),
    .Y(_08300_));
 sky130_fd_sc_hd__o21a_2 _36248_ (.A1(_08298_),
    .A2(_08299_),
    .B1(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__nor3_2 _36249_ (.A(_08298_),
    .B(_08299_),
    .C(_08300_),
    .Y(_08302_));
 sky130_fd_sc_hd__nor2_2 _36250_ (.A(_08301_),
    .B(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__o21ai_2 _36251_ (.A1(_08056_),
    .A2(_08060_),
    .B1(_08303_),
    .Y(_08304_));
 sky130_fd_sc_hd__or3_2 _36252_ (.A(_08056_),
    .B(_08060_),
    .C(_08303_),
    .X(_08305_));
 sky130_fd_sc_hd__and2_2 _36253_ (.A(_08304_),
    .B(_08305_),
    .X(_08307_));
 sky130_fd_sc_hd__xnor2_2 _36254_ (.A(_08297_),
    .B(_08307_),
    .Y(_08308_));
 sky130_fd_sc_hd__o21a_2 _36255_ (.A1(_08070_),
    .A2(_08073_),
    .B1(_08308_),
    .X(_08309_));
 sky130_fd_sc_hd__nor3_2 _36256_ (.A(_08070_),
    .B(_08073_),
    .C(_08308_),
    .Y(_08310_));
 sky130_fd_sc_hd__a211oi_2 _36257_ (.A1(_08294_),
    .A2(_08296_),
    .B1(_08309_),
    .C1(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__o211a_2 _36258_ (.A1(_08309_),
    .A2(_08310_),
    .B1(_08294_),
    .C1(_08296_),
    .X(_08312_));
 sky130_fd_sc_hd__nor2_2 _36259_ (.A(_08114_),
    .B(_08116_),
    .Y(_08313_));
 sky130_fd_sc_hd__or3_2 _36260_ (.A(_08311_),
    .B(_08312_),
    .C(_08313_),
    .X(_08314_));
 sky130_fd_sc_hd__o21ai_2 _36261_ (.A1(_08311_),
    .A2(_08312_),
    .B1(_08313_),
    .Y(_08315_));
 sky130_fd_sc_hd__nand3_2 _36262_ (.A(_08293_),
    .B(_08314_),
    .C(_08315_),
    .Y(_08316_));
 sky130_fd_sc_hd__a21o_2 _36263_ (.A1(_08314_),
    .A2(_08315_),
    .B1(_08293_),
    .X(_08318_));
 sky130_fd_sc_hd__and3_2 _36264_ (.A(_08080_),
    .B(_08316_),
    .C(_08318_),
    .X(_08319_));
 sky130_fd_sc_hd__a21oi_2 _36265_ (.A1(_08316_),
    .A2(_08318_),
    .B1(_08080_),
    .Y(_08320_));
 sky130_fd_sc_hd__a211oi_2 _36266_ (.A1(_08119_),
    .A2(_08272_),
    .B1(_08319_),
    .C1(_08320_),
    .Y(_08321_));
 sky130_fd_sc_hd__o211a_2 _36267_ (.A1(_08319_),
    .A2(_08320_),
    .B1(_08119_),
    .C1(_08272_),
    .X(_08322_));
 sky130_fd_sc_hd__nor3_2 _36268_ (.A(_08271_),
    .B(_08321_),
    .C(_08322_),
    .Y(_08323_));
 sky130_fd_sc_hd__o21a_2 _36269_ (.A1(_08321_),
    .A2(_08322_),
    .B1(_08271_),
    .X(_08324_));
 sky130_fd_sc_hd__or3_2 _36270_ (.A(_08129_),
    .B(_08323_),
    .C(_08324_),
    .X(_08325_));
 sky130_fd_sc_hd__o21ai_2 _36271_ (.A1(_08323_),
    .A2(_08324_),
    .B1(_08129_),
    .Y(_08326_));
 sky130_fd_sc_hd__o211ai_2 _36272_ (.A1(_08124_),
    .A2(_08127_),
    .B1(_08325_),
    .C1(_08326_),
    .Y(_08327_));
 sky130_fd_sc_hd__a211o_2 _36273_ (.A1(_08325_),
    .A2(_08326_),
    .B1(_08124_),
    .C1(_08127_),
    .X(_08329_));
 sky130_fd_sc_hd__and2_2 _36274_ (.A(_08327_),
    .B(_08329_),
    .X(_08330_));
 sky130_fd_sc_hd__or2_2 _36275_ (.A(_08132_),
    .B(_08134_),
    .X(_08331_));
 sky130_fd_sc_hd__xnor2_2 _36276_ (.A(_08330_),
    .B(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__o21ba_2 _36277_ (.A1(_08094_),
    .A2(_08099_),
    .B1_N(_08332_),
    .X(_08333_));
 sky130_fd_sc_hd__or3b_2 _36278_ (.A(_08094_),
    .B(_08099_),
    .C_N(_08332_),
    .X(_08334_));
 sky130_fd_sc_hd__or2b_2 _36279_ (.A(_08333_),
    .B_N(_08334_),
    .X(_08335_));
 sky130_fd_sc_hd__nor2_2 _36280_ (.A(_08136_),
    .B(_08138_),
    .Y(_08336_));
 sky130_fd_sc_hd__nor2_2 _36281_ (.A(_08335_),
    .B(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__and2_2 _36282_ (.A(_08335_),
    .B(_08336_),
    .X(_08338_));
 sky130_fd_sc_hd__nor2_2 _36283_ (.A(_08337_),
    .B(_08338_),
    .Y(_08340_));
 sky130_fd_sc_hd__o21bai_2 _36284_ (.A1(_07903_),
    .A2(_08141_),
    .B1_N(_08143_),
    .Y(_08341_));
 sky130_fd_sc_hd__o31a_2 _36285_ (.A1(_07905_),
    .A2(_07910_),
    .A3(_08144_),
    .B1(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__xor2_2 _36286_ (.A(_08340_),
    .B(_08342_),
    .X(_08343_));
 sky130_fd_sc_hd__and3_2 _36287_ (.A(_08253_),
    .B(_08254_),
    .C(_08343_),
    .X(_08344_));
 sky130_fd_sc_hd__a21oi_2 _36288_ (.A1(_08253_),
    .A2(_08254_),
    .B1(_08343_),
    .Y(_08345_));
 sky130_fd_sc_hd__nor2_2 _36289_ (.A(_08344_),
    .B(_08345_),
    .Y(_08346_));
 sky130_fd_sc_hd__xor2_2 _36290_ (.A(_16226_),
    .B(_08346_),
    .X(_08347_));
 sky130_fd_sc_hd__nand2_2 _36291_ (.A(_16134_),
    .B(_08147_),
    .Y(_08348_));
 sky130_fd_sc_hd__o21a_2 _36292_ (.A1(_08053_),
    .A2(_08146_),
    .B1(_08348_),
    .X(_08349_));
 sky130_fd_sc_hd__nor2_2 _36293_ (.A(_08347_),
    .B(_08349_),
    .Y(_08351_));
 sky130_fd_sc_hd__and2_2 _36294_ (.A(_08347_),
    .B(_08349_),
    .X(_08352_));
 sky130_fd_sc_hd__or2_2 _36295_ (.A(_08351_),
    .B(_08352_),
    .X(_08353_));
 sky130_fd_sc_hd__nand2_2 _36296_ (.A(_07918_),
    .B(_08151_),
    .Y(_08354_));
 sky130_fd_sc_hd__a31o_2 _36297_ (.A1(_07921_),
    .A2(_07923_),
    .A3(_07927_),
    .B1(_08354_),
    .X(_08355_));
 sky130_fd_sc_hd__nand2_2 _36298_ (.A(_08148_),
    .B(_08150_),
    .Y(_08356_));
 sky130_fd_sc_hd__nor2_2 _36299_ (.A(_08148_),
    .B(_08150_),
    .Y(_08357_));
 sky130_fd_sc_hd__a21oi_2 _36300_ (.A1(_07916_),
    .A2(_08356_),
    .B1(_08357_),
    .Y(_08358_));
 sky130_fd_sc_hd__and2_2 _36301_ (.A(_08355_),
    .B(_08358_),
    .X(_08359_));
 sky130_fd_sc_hd__xor2_2 _36302_ (.A(_08353_),
    .B(_08359_),
    .X(_08360_));
 sky130_fd_sc_hd__xnor2_2 _36303_ (.A(_16463_),
    .B(_08360_),
    .Y(_08362_));
 sky130_fd_sc_hd__a21oi_2 _36304_ (.A1(_07930_),
    .A2(_08157_),
    .B1(_08156_),
    .Y(_08363_));
 sky130_fd_sc_hd__a21o_2 _36305_ (.A1(_07947_),
    .A2(_08158_),
    .B1(_08363_),
    .X(_08364_));
 sky130_fd_sc_hd__xor2_2 _36306_ (.A(_08362_),
    .B(_08364_),
    .X(oO[82]));
 sky130_fd_sc_hd__o21bai_2 _36307_ (.A1(_08353_),
    .A2(_08359_),
    .B1_N(_08351_),
    .Y(_08365_));
 sky130_fd_sc_hd__or2_2 _36308_ (.A(_08248_),
    .B(_08250_),
    .X(_08366_));
 sky130_fd_sc_hd__or2b_2 _36309_ (.A(_08246_),
    .B_N(_08245_),
    .X(_08367_));
 sky130_fd_sc_hd__nand2_2 _36310_ (.A(_08160_),
    .B(_08247_),
    .Y(_08368_));
 sky130_fd_sc_hd__o21a_2 _36311_ (.A1(_08241_),
    .A2(_08242_),
    .B1(_08239_),
    .X(_08369_));
 sky130_fd_sc_hd__or2b_2 _36312_ (.A(_08235_),
    .B_N(_08237_),
    .X(_08370_));
 sky130_fd_sc_hd__nand2_2 _36313_ (.A(_08238_),
    .B(_08244_),
    .Y(_08372_));
 sky130_fd_sc_hd__or2_2 _36314_ (.A(_08161_),
    .B(_08178_),
    .X(_08373_));
 sky130_fd_sc_hd__or2_2 _36315_ (.A(_08179_),
    .B(_08234_),
    .X(_08374_));
 sky130_fd_sc_hd__and3_2 _36316_ (.A(_08167_),
    .B(_08168_),
    .C(_08177_),
    .X(_08375_));
 sky130_fd_sc_hd__and4_2 _36317_ (.A(_06414_),
    .B(_06411_),
    .C(_03458_),
    .D(_04905_),
    .X(_08376_));
 sky130_fd_sc_hd__o22a_2 _36318_ (.A1(_05978_),
    .A2(_06797_),
    .B1(_05550_),
    .B2(_05980_),
    .X(_08377_));
 sky130_fd_sc_hd__nor2_2 _36319_ (.A(_08376_),
    .B(_08377_),
    .Y(_08378_));
 sky130_fd_sc_hd__nand2_2 _36320_ (.A(_06813_),
    .B(_06154_),
    .Y(_08379_));
 sky130_fd_sc_hd__xnor2_2 _36321_ (.A(_08378_),
    .B(_08379_),
    .Y(_08380_));
 sky130_fd_sc_hd__nand2_2 _36322_ (.A(_05533_),
    .B(_03938_),
    .Y(_08381_));
 sky130_fd_sc_hd__o22a_2 _36323_ (.A1(_05983_),
    .A2(_06786_),
    .B1(_08164_),
    .B2(_04847_),
    .X(_08383_));
 sky130_fd_sc_hd__a21o_2 _36324_ (.A1(_05533_),
    .A2(_04844_),
    .B1(_08383_),
    .X(_08384_));
 sky130_fd_sc_hd__a21o_2 _36325_ (.A1(_08381_),
    .A2(_08167_),
    .B1(_08384_),
    .X(_08385_));
 sky130_fd_sc_hd__nand3_2 _36326_ (.A(_08381_),
    .B(_08167_),
    .C(_08384_),
    .Y(_08386_));
 sky130_fd_sc_hd__nand3_2 _36327_ (.A(_08380_),
    .B(_08385_),
    .C(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__a21o_2 _36328_ (.A1(_08385_),
    .A2(_08386_),
    .B1(_08380_),
    .X(_08388_));
 sky130_fd_sc_hd__nand3_2 _36329_ (.A(_08375_),
    .B(_08387_),
    .C(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__a21o_2 _36330_ (.A1(_08387_),
    .A2(_08388_),
    .B1(_08375_),
    .X(_08390_));
 sky130_fd_sc_hd__and2b_2 _36331_ (.A_N(_08215_),
    .B(_08209_),
    .X(_08391_));
 sky130_fd_sc_hd__and2b_2 _36332_ (.A_N(_08208_),
    .B(_08216_),
    .X(_08392_));
 sky130_fd_sc_hd__buf_1 _36333_ (.A(_05550_),
    .X(_08394_));
 sky130_fd_sc_hd__a211o_2 _36334_ (.A1(_07468_),
    .A2(_08175_),
    .B1(_04847_),
    .C1(_08394_),
    .X(_08395_));
 sky130_fd_sc_hd__a21bo_2 _36335_ (.A1(_08212_),
    .A2(_08214_),
    .B1_N(_08211_),
    .X(_08396_));
 sky130_fd_sc_hd__nand2_2 _36336_ (.A(_07039_),
    .B(_07472_),
    .Y(_08397_));
 sky130_fd_sc_hd__xor2_2 _36337_ (.A(_08210_),
    .B(_08397_),
    .X(_08398_));
 sky130_fd_sc_hd__nand2_2 _36338_ (.A(_06484_),
    .B(_06983_),
    .Y(_08399_));
 sky130_fd_sc_hd__xor2_2 _36339_ (.A(_08398_),
    .B(_08399_),
    .X(_08400_));
 sky130_fd_sc_hd__a21bo_2 _36340_ (.A1(_08171_),
    .A2(_08173_),
    .B1_N(_08170_),
    .X(_08401_));
 sky130_fd_sc_hd__and2b_2 _36341_ (.A_N(_08400_),
    .B(_08401_),
    .X(_08402_));
 sky130_fd_sc_hd__and2b_2 _36342_ (.A_N(_08401_),
    .B(_08400_),
    .X(_08403_));
 sky130_fd_sc_hd__nor2_2 _36343_ (.A(_08402_),
    .B(_08403_),
    .Y(_08405_));
 sky130_fd_sc_hd__xnor2_2 _36344_ (.A(_08396_),
    .B(_08405_),
    .Y(_08406_));
 sky130_fd_sc_hd__xor2_2 _36345_ (.A(_08395_),
    .B(_08406_),
    .X(_08407_));
 sky130_fd_sc_hd__o21ai_2 _36346_ (.A1(_08391_),
    .A2(_08392_),
    .B1(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__or3_2 _36347_ (.A(_08391_),
    .B(_08392_),
    .C(_08407_),
    .X(_08409_));
 sky130_fd_sc_hd__nand2_2 _36348_ (.A(_08408_),
    .B(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__a21o_2 _36349_ (.A1(_08219_),
    .A2(_08222_),
    .B1(_08410_),
    .X(_08411_));
 sky130_fd_sc_hd__nand3_2 _36350_ (.A(_08219_),
    .B(_08222_),
    .C(_08410_),
    .Y(_08412_));
 sky130_fd_sc_hd__nand2_2 _36351_ (.A(_08411_),
    .B(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__a21o_2 _36352_ (.A1(_08184_),
    .A2(_08186_),
    .B1(_08182_),
    .X(_08414_));
 sky130_fd_sc_hd__nor2_2 _36353_ (.A(_04862_),
    .B(_05931_),
    .Y(_08416_));
 sky130_fd_sc_hd__and3_2 _36354_ (.A(_05507_),
    .B(_04781_),
    .C(_08416_),
    .X(_08417_));
 sky130_fd_sc_hd__o22a_2 _36355_ (.A1(_04862_),
    .A2(_04782_),
    .B1(_07252_),
    .B2(_05979_),
    .X(_08418_));
 sky130_fd_sc_hd__nor2_2 _36356_ (.A(_08417_),
    .B(_08418_),
    .Y(_08419_));
 sky130_fd_sc_hd__nor2_2 _36357_ (.A(_04501_),
    .B(_05440_),
    .Y(_08420_));
 sky130_fd_sc_hd__xor2_2 _36358_ (.A(_08419_),
    .B(_08420_),
    .X(_08421_));
 sky130_fd_sc_hd__nand2_2 _36359_ (.A(_06822_),
    .B(_05450_),
    .Y(_08422_));
 sky130_fd_sc_hd__xnor2_2 _36360_ (.A(_08188_),
    .B(_08422_),
    .Y(_08423_));
 sky130_fd_sc_hd__or3_2 _36361_ (.A(_05504_),
    .B(_00944_),
    .C(_08423_),
    .X(_08424_));
 sky130_fd_sc_hd__o21ai_2 _36362_ (.A1(_05504_),
    .A2(_00944_),
    .B1(_08423_),
    .Y(_08425_));
 sky130_fd_sc_hd__nand2_2 _36363_ (.A(_08424_),
    .B(_08425_),
    .Y(_08427_));
 sky130_fd_sc_hd__o22a_2 _36364_ (.A1(_07992_),
    .A2(_08188_),
    .B1(_08189_),
    .B2(_08191_),
    .X(_08428_));
 sky130_fd_sc_hd__or2_2 _36365_ (.A(_08427_),
    .B(_08428_),
    .X(_08429_));
 sky130_fd_sc_hd__nand2_2 _36366_ (.A(_08427_),
    .B(_08428_),
    .Y(_08430_));
 sky130_fd_sc_hd__and2_2 _36367_ (.A(_08429_),
    .B(_08430_),
    .X(_08431_));
 sky130_fd_sc_hd__nand2_2 _36368_ (.A(_08421_),
    .B(_08431_),
    .Y(_08432_));
 sky130_fd_sc_hd__or2_2 _36369_ (.A(_08421_),
    .B(_08431_),
    .X(_08433_));
 sky130_fd_sc_hd__nand2_2 _36370_ (.A(_08432_),
    .B(_08433_),
    .Y(_08434_));
 sky130_fd_sc_hd__a21oi_2 _36371_ (.A1(_08194_),
    .A2(_08198_),
    .B1(_08434_),
    .Y(_08435_));
 sky130_fd_sc_hd__and3_2 _36372_ (.A(_08194_),
    .B(_08198_),
    .C(_08434_),
    .X(_08436_));
 sky130_fd_sc_hd__nor2_2 _36373_ (.A(_08435_),
    .B(_08436_),
    .Y(_08438_));
 sky130_fd_sc_hd__xnor2_2 _36374_ (.A(_08414_),
    .B(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__xnor2_2 _36375_ (.A(_08413_),
    .B(_08439_),
    .Y(_08440_));
 sky130_fd_sc_hd__a21oi_2 _36376_ (.A1(_08225_),
    .A2(_08227_),
    .B1(_08440_),
    .Y(_08441_));
 sky130_fd_sc_hd__and3_2 _36377_ (.A(_08225_),
    .B(_08227_),
    .C(_08440_),
    .X(_08442_));
 sky130_fd_sc_hd__nor2_2 _36378_ (.A(_08441_),
    .B(_08442_),
    .Y(_08443_));
 sky130_fd_sc_hd__and3_2 _36379_ (.A(_08389_),
    .B(_08390_),
    .C(_08443_),
    .X(_08444_));
 sky130_fd_sc_hd__a21oi_2 _36380_ (.A1(_08389_),
    .A2(_08390_),
    .B1(_08443_),
    .Y(_08445_));
 sky130_fd_sc_hd__a211o_2 _36381_ (.A1(_08373_),
    .A2(_08374_),
    .B1(_08444_),
    .C1(_08445_),
    .X(_08446_));
 sky130_fd_sc_hd__o211ai_2 _36382_ (.A1(_08444_),
    .A2(_08445_),
    .B1(_08373_),
    .C1(_08374_),
    .Y(_08447_));
 sky130_fd_sc_hd__or2_2 _36383_ (.A(_08230_),
    .B(_08232_),
    .X(_08449_));
 sky130_fd_sc_hd__and3_2 _36384_ (.A(_08198_),
    .B(_08199_),
    .C(_08201_),
    .X(_08450_));
 sky130_fd_sc_hd__and2b_2 _36385_ (.A_N(_08180_),
    .B(_08202_),
    .X(_08451_));
 sky130_fd_sc_hd__nor2_2 _36386_ (.A(_08450_),
    .B(_08451_),
    .Y(_08452_));
 sky130_fd_sc_hd__xnor2_2 _36387_ (.A(_08449_),
    .B(_08452_),
    .Y(_08453_));
 sky130_fd_sc_hd__and3_2 _36388_ (.A(_08446_),
    .B(_08447_),
    .C(_08453_),
    .X(_08454_));
 sky130_fd_sc_hd__a21oi_2 _36389_ (.A1(_08446_),
    .A2(_08447_),
    .B1(_08453_),
    .Y(_08455_));
 sky130_fd_sc_hd__a211o_2 _36390_ (.A1(_08370_),
    .A2(_08372_),
    .B1(_08454_),
    .C1(_08455_),
    .X(_08456_));
 sky130_fd_sc_hd__o211ai_2 _36391_ (.A1(_08454_),
    .A2(_08455_),
    .B1(_08370_),
    .C1(_08372_),
    .Y(_08457_));
 sky130_fd_sc_hd__and3_2 _36392_ (.A(_08369_),
    .B(_08456_),
    .C(_08457_),
    .X(_08458_));
 sky130_fd_sc_hd__a21oi_2 _36393_ (.A1(_08456_),
    .A2(_08457_),
    .B1(_08369_),
    .Y(_08460_));
 sky130_fd_sc_hd__a211oi_2 _36394_ (.A1(_08367_),
    .A2(_08368_),
    .B1(_08458_),
    .C1(_08460_),
    .Y(_08461_));
 sky130_fd_sc_hd__o211a_2 _36395_ (.A1(_08458_),
    .A2(_08460_),
    .B1(_08367_),
    .C1(_08368_),
    .X(_08462_));
 sky130_fd_sc_hd__nor2_2 _36396_ (.A(_08461_),
    .B(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__nand3_2 _36397_ (.A(_08366_),
    .B(_08253_),
    .C(_08463_),
    .Y(_08464_));
 sky130_fd_sc_hd__a21o_2 _36398_ (.A1(_08366_),
    .A2(_08253_),
    .B1(_08463_),
    .X(_08465_));
 sky130_fd_sc_hd__and2_2 _36399_ (.A(_08330_),
    .B(_08331_),
    .X(_08466_));
 sky130_fd_sc_hd__and3b_2 _36400_ (.A_N(_07820_),
    .B(iX[63]),
    .C(iY[52]),
    .X(_08467_));
 sky130_fd_sc_hd__and2_2 _36401_ (.A(iY[54]),
    .B(iX[62]),
    .X(_08468_));
 sky130_fd_sc_hd__and3_2 _36402_ (.A(iY[53]),
    .B(iX[61]),
    .C(_08468_),
    .X(_08469_));
 sky130_fd_sc_hd__a22oi_2 _36403_ (.A1(iY[54]),
    .A2(iX[61]),
    .B1(iX[62]),
    .B2(iY[53]),
    .Y(_08471_));
 sky130_fd_sc_hd__nor2_2 _36404_ (.A(_08469_),
    .B(_08471_),
    .Y(_08472_));
 sky130_fd_sc_hd__a21oi_2 _36405_ (.A1(iY[55]),
    .A2(iX[60]),
    .B1(_08472_),
    .Y(_08473_));
 sky130_fd_sc_hd__and3_2 _36406_ (.A(iY[55]),
    .B(iX[60]),
    .C(_08472_),
    .X(_08474_));
 sky130_fd_sc_hd__nor2_2 _36407_ (.A(_08473_),
    .B(_08474_),
    .Y(_08475_));
 sky130_fd_sc_hd__xnor2_2 _36408_ (.A(_08467_),
    .B(_08475_),
    .Y(_08476_));
 sky130_fd_sc_hd__or2b_2 _36409_ (.A(_08279_),
    .B_N(_08278_),
    .X(_08477_));
 sky130_fd_sc_hd__and4_2 _36410_ (.A(iX[55]),
    .B(iX[56]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_08478_));
 sky130_fd_sc_hd__a22oi_2 _36411_ (.A1(iX[56]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[55]),
    .Y(_08479_));
 sky130_fd_sc_hd__nor2_2 _36412_ (.A(_08478_),
    .B(_08479_),
    .Y(_08480_));
 sky130_fd_sc_hd__nand2_2 _36413_ (.A(iX[54]),
    .B(iY[61]),
    .Y(_08482_));
 sky130_fd_sc_hd__xnor2_2 _36414_ (.A(_08480_),
    .B(_08482_),
    .Y(_08483_));
 sky130_fd_sc_hd__o21ba_2 _36415_ (.A1(_08275_),
    .A2(_08277_),
    .B1_N(_08274_),
    .X(_08484_));
 sky130_fd_sc_hd__xnor2_2 _36416_ (.A(_08483_),
    .B(_08484_),
    .Y(_08485_));
 sky130_fd_sc_hd__and2_2 _36417_ (.A(iX[53]),
    .B(iY[62]),
    .X(_08486_));
 sky130_fd_sc_hd__or2_2 _36418_ (.A(_08485_),
    .B(_08486_),
    .X(_08487_));
 sky130_fd_sc_hd__nand2_2 _36419_ (.A(_08485_),
    .B(_08486_),
    .Y(_08488_));
 sky130_fd_sc_hd__nand2_2 _36420_ (.A(_08487_),
    .B(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__a21oi_2 _36421_ (.A1(_08477_),
    .A2(_08283_),
    .B1(_08489_),
    .Y(_08490_));
 sky130_fd_sc_hd__and3_2 _36422_ (.A(_08477_),
    .B(_08283_),
    .C(_08489_),
    .X(_08491_));
 sky130_fd_sc_hd__nor2_2 _36423_ (.A(_08490_),
    .B(_08491_),
    .Y(_08493_));
 sky130_fd_sc_hd__nand2_2 _36424_ (.A(iX[52]),
    .B(iY[63]),
    .Y(_08494_));
 sky130_fd_sc_hd__xnor2_2 _36425_ (.A(_08493_),
    .B(_08494_),
    .Y(_08495_));
 sky130_fd_sc_hd__or2b_2 _36426_ (.A(_08297_),
    .B_N(_08307_),
    .X(_08496_));
 sky130_fd_sc_hd__or2b_2 _36427_ (.A(_08257_),
    .B_N(_08258_),
    .X(_08497_));
 sky130_fd_sc_hd__o21ba_2 _36428_ (.A1(_08261_),
    .A2(_08264_),
    .B1_N(_08260_),
    .X(_08498_));
 sky130_fd_sc_hd__and4_2 _36429_ (.A(iY[56]),
    .B(iY[57]),
    .C(iX[58]),
    .D(iX[59]),
    .X(_08499_));
 sky130_fd_sc_hd__a22oi_2 _36430_ (.A1(iY[57]),
    .A2(iX[58]),
    .B1(iX[59]),
    .B2(iY[56]),
    .Y(_08500_));
 sky130_fd_sc_hd__nor2_2 _36431_ (.A(_08499_),
    .B(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__nand2_2 _36432_ (.A(iX[57]),
    .B(iY[58]),
    .Y(_08502_));
 sky130_fd_sc_hd__xnor2_2 _36433_ (.A(_08501_),
    .B(_08502_),
    .Y(_08504_));
 sky130_fd_sc_hd__xnor2_2 _36434_ (.A(_08498_),
    .B(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__o21a_2 _36435_ (.A1(_08298_),
    .A2(_08302_),
    .B1(_08505_),
    .X(_08506_));
 sky130_fd_sc_hd__nor3_2 _36436_ (.A(_08298_),
    .B(_08302_),
    .C(_08505_),
    .Y(_08507_));
 sky130_fd_sc_hd__or2_2 _36437_ (.A(_08506_),
    .B(_08507_),
    .X(_08508_));
 sky130_fd_sc_hd__a21oi_2 _36438_ (.A1(_08497_),
    .A2(_08266_),
    .B1(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__and3_2 _36439_ (.A(_08497_),
    .B(_08266_),
    .C(_08508_),
    .X(_08510_));
 sky130_fd_sc_hd__a211o_2 _36440_ (.A1(_08304_),
    .A2(_08496_),
    .B1(_08509_),
    .C1(_08510_),
    .X(_08511_));
 sky130_fd_sc_hd__o211ai_2 _36441_ (.A1(_08509_),
    .A2(_08510_),
    .B1(_08304_),
    .C1(_08496_),
    .Y(_08512_));
 sky130_fd_sc_hd__o211ai_2 _36442_ (.A1(_08309_),
    .A2(_08311_),
    .B1(_08511_),
    .C1(_08512_),
    .Y(_08513_));
 sky130_fd_sc_hd__a211o_2 _36443_ (.A1(_08511_),
    .A2(_08512_),
    .B1(_08309_),
    .C1(_08311_),
    .X(_08515_));
 sky130_fd_sc_hd__and3_2 _36444_ (.A(_08495_),
    .B(_08513_),
    .C(_08515_),
    .X(_08516_));
 sky130_fd_sc_hd__a21oi_2 _36445_ (.A1(_08513_),
    .A2(_08515_),
    .B1(_08495_),
    .Y(_08517_));
 sky130_fd_sc_hd__nor3_2 _36446_ (.A(_08269_),
    .B(_08516_),
    .C(_08517_),
    .Y(_08518_));
 sky130_fd_sc_hd__o21a_2 _36447_ (.A1(_08516_),
    .A2(_08517_),
    .B1(_08269_),
    .X(_08519_));
 sky130_fd_sc_hd__a211oi_2 _36448_ (.A1(_08314_),
    .A2(_08316_),
    .B1(_08518_),
    .C1(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__o211a_2 _36449_ (.A1(_08518_),
    .A2(_08519_),
    .B1(_08314_),
    .C1(_08316_),
    .X(_08521_));
 sky130_fd_sc_hd__or3_2 _36450_ (.A(_08476_),
    .B(_08520_),
    .C(_08521_),
    .X(_08522_));
 sky130_fd_sc_hd__o21ai_2 _36451_ (.A1(_08520_),
    .A2(_08521_),
    .B1(_08476_),
    .Y(_08523_));
 sky130_fd_sc_hd__and3_2 _36452_ (.A(_08323_),
    .B(_08522_),
    .C(_08523_),
    .X(_08524_));
 sky130_fd_sc_hd__a21oi_2 _36453_ (.A1(_08522_),
    .A2(_08523_),
    .B1(_08323_),
    .Y(_08526_));
 sky130_fd_sc_hd__nor2_2 _36454_ (.A(_08524_),
    .B(_08526_),
    .Y(_08527_));
 sky130_fd_sc_hd__o21a_2 _36455_ (.A1(_08319_),
    .A2(_08321_),
    .B1(_08527_),
    .X(_08528_));
 sky130_fd_sc_hd__nor3_2 _36456_ (.A(_08319_),
    .B(_08321_),
    .C(_08527_),
    .Y(_08529_));
 sky130_fd_sc_hd__a211oi_2 _36457_ (.A1(_08325_),
    .A2(_08327_),
    .B1(_08528_),
    .C1(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__o211a_2 _36458_ (.A1(_08528_),
    .A2(_08529_),
    .B1(_08325_),
    .C1(_08327_),
    .X(_08531_));
 sky130_fd_sc_hd__a211oi_2 _36459_ (.A1(_08287_),
    .A2(_08292_),
    .B1(_08530_),
    .C1(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__o211a_2 _36460_ (.A1(_08530_),
    .A2(_08531_),
    .B1(_08287_),
    .C1(_08292_),
    .X(_08533_));
 sky130_fd_sc_hd__nor2_2 _36461_ (.A(_08532_),
    .B(_08533_),
    .Y(_08534_));
 sky130_fd_sc_hd__or3_2 _36462_ (.A(_08466_),
    .B(_08333_),
    .C(_08534_),
    .X(_08535_));
 sky130_fd_sc_hd__o21ai_2 _36463_ (.A1(_08466_),
    .A2(_08333_),
    .B1(_08534_),
    .Y(_08537_));
 sky130_fd_sc_hd__and2_2 _36464_ (.A(_08535_),
    .B(_08537_),
    .X(_08538_));
 sky130_fd_sc_hd__o21ba_2 _36465_ (.A1(_08338_),
    .A2(_08342_),
    .B1_N(_08337_),
    .X(_08539_));
 sky130_fd_sc_hd__xnor2_2 _36466_ (.A(_08538_),
    .B(_08539_),
    .Y(_08540_));
 sky130_fd_sc_hd__nand3_2 _36467_ (.A(_08464_),
    .B(_08465_),
    .C(_08540_),
    .Y(_08541_));
 sky130_fd_sc_hd__a21o_2 _36468_ (.A1(_08464_),
    .A2(_08465_),
    .B1(_08540_),
    .X(_08542_));
 sky130_fd_sc_hd__nand3_2 _36469_ (.A(_16809_),
    .B(_08541_),
    .C(_08542_),
    .Y(_08543_));
 sky130_fd_sc_hd__a21o_2 _36470_ (.A1(_08541_),
    .A2(_08542_),
    .B1(_16809_),
    .X(_08544_));
 sky130_fd_sc_hd__o21bai_2 _36471_ (.A1(_16226_),
    .A2(_08345_),
    .B1_N(_08344_),
    .Y(_08545_));
 sky130_fd_sc_hd__a21oi_2 _36472_ (.A1(_08543_),
    .A2(_08544_),
    .B1(_08545_),
    .Y(_08546_));
 sky130_fd_sc_hd__nand3_2 _36473_ (.A(_08545_),
    .B(_08543_),
    .C(_08544_),
    .Y(_08548_));
 sky130_fd_sc_hd__and2b_2 _36474_ (.A_N(_08546_),
    .B(_08548_),
    .X(_08549_));
 sky130_fd_sc_hd__xnor2_2 _36475_ (.A(_08365_),
    .B(_08549_),
    .Y(_08550_));
 sky130_fd_sc_hd__nor2_2 _36476_ (.A(_16597_),
    .B(_08550_),
    .Y(_08551_));
 sky130_fd_sc_hd__nand2_2 _36477_ (.A(_16597_),
    .B(_08550_),
    .Y(_08552_));
 sky130_fd_sc_hd__and2b_2 _36478_ (.A_N(_08551_),
    .B(_08552_),
    .X(_08553_));
 sky130_fd_sc_hd__and2b_2 _36479_ (.A_N(_16463_),
    .B(_08360_),
    .X(_08554_));
 sky130_fd_sc_hd__a21oi_2 _36480_ (.A1(_08362_),
    .A2(_08364_),
    .B1(_08554_),
    .Y(_08555_));
 sky130_fd_sc_hd__xnor2_2 _36481_ (.A(_08553_),
    .B(_08555_),
    .Y(oO[83]));
 sky130_fd_sc_hd__and2_2 _36482_ (.A(_08362_),
    .B(_08553_),
    .X(_08556_));
 sky130_fd_sc_hd__a21oi_2 _36483_ (.A1(_08554_),
    .A2(_08552_),
    .B1(_08551_),
    .Y(_08558_));
 sky130_fd_sc_hd__a21boi_2 _36484_ (.A1(_08364_),
    .A2(_08556_),
    .B1_N(_08558_),
    .Y(_08559_));
 sky130_fd_sc_hd__o21a_2 _36485_ (.A1(_08450_),
    .A2(_08451_),
    .B1(_08449_),
    .X(_08560_));
 sky130_fd_sc_hd__or2_2 _36486_ (.A(_06399_),
    .B(_05495_),
    .X(_08561_));
 sky130_fd_sc_hd__a2bb2o_2 _36487_ (.A1_N(_04501_),
    .A2_N(_06786_),
    .B1(_04005_),
    .B2(_06414_),
    .X(_08562_));
 sky130_fd_sc_hd__nand2_2 _36488_ (.A(_08561_),
    .B(_08562_),
    .Y(_08563_));
 sky130_fd_sc_hd__inv_2 _36489_ (.A(_08384_),
    .Y(_08564_));
 sky130_fd_sc_hd__inv_2 _36490_ (.A(_08162_),
    .Y(_08565_));
 sky130_fd_sc_hd__o2bb2a_2 _36491_ (.A1_N(_05533_),
    .A2_N(_04844_),
    .B1(_08165_),
    .B2(_08565_),
    .X(_08566_));
 sky130_fd_sc_hd__a21oi_2 _36492_ (.A1(_08381_),
    .A2(_08566_),
    .B1(_08383_),
    .Y(_08567_));
 sky130_fd_sc_hd__a31o_2 _36493_ (.A1(_07975_),
    .A2(_08166_),
    .A3(_08564_),
    .B1(_08567_),
    .X(_08569_));
 sky130_fd_sc_hd__xor2_2 _36494_ (.A(_08563_),
    .B(_08569_),
    .X(_08570_));
 sky130_fd_sc_hd__buf_1 _36495_ (.A(_06797_),
    .X(_08571_));
 sky130_fd_sc_hd__o22a_2 _36496_ (.A1(_05500_),
    .A2(_08571_),
    .B1(_08394_),
    .B2(_05978_),
    .X(_08572_));
 sky130_fd_sc_hd__and4_2 _36497_ (.A(_06411_),
    .B(_06813_),
    .C(_03458_),
    .D(_04905_),
    .X(_08573_));
 sky130_fd_sc_hd__or2_2 _36498_ (.A(_08572_),
    .B(_08573_),
    .X(_08574_));
 sky130_fd_sc_hd__xor2_2 _36499_ (.A(_08570_),
    .B(_08574_),
    .X(_08575_));
 sky130_fd_sc_hd__xnor2_2 _36500_ (.A(_08387_),
    .B(_08575_),
    .Y(_08576_));
 sky130_fd_sc_hd__or3b_2 _36501_ (.A(_03341_),
    .B(_05227_),
    .C_N(_08398_),
    .X(_08577_));
 sky130_fd_sc_hd__o21a_2 _36502_ (.A1(_08210_),
    .A2(_08397_),
    .B1(_08577_),
    .X(_08578_));
 sky130_fd_sc_hd__o21ba_2 _36503_ (.A1(_08377_),
    .A2(_08379_),
    .B1_N(_08376_),
    .X(_08580_));
 sky130_fd_sc_hd__and4_2 _36504_ (.A(_07039_),
    .B(_06488_),
    .C(_07472_),
    .D(_06154_),
    .X(_08581_));
 sky130_fd_sc_hd__buf_1 _36505_ (.A(_05231_),
    .X(_08582_));
 sky130_fd_sc_hd__o22a_2 _36506_ (.A1(_18344_),
    .A2(_06023_),
    .B1(_08582_),
    .B2(_06491_),
    .X(_08583_));
 sky130_fd_sc_hd__nor2_2 _36507_ (.A(_08581_),
    .B(_08583_),
    .Y(_08584_));
 sky130_fd_sc_hd__and3_2 _36508_ (.A(_07279_),
    .B(_07461_),
    .C(_08584_),
    .X(_08585_));
 sky130_fd_sc_hd__a21oi_2 _36509_ (.A1(_07279_),
    .A2(_07461_),
    .B1(_08584_),
    .Y(_08586_));
 sky130_fd_sc_hd__nor2_2 _36510_ (.A(_08585_),
    .B(_08586_),
    .Y(_08587_));
 sky130_fd_sc_hd__xnor2_2 _36511_ (.A(_08580_),
    .B(_08587_),
    .Y(_08588_));
 sky130_fd_sc_hd__or2b_2 _36512_ (.A(_08578_),
    .B_N(_08588_),
    .X(_08589_));
 sky130_fd_sc_hd__or2b_2 _36513_ (.A(_08588_),
    .B_N(_08578_),
    .X(_08591_));
 sky130_fd_sc_hd__nand2_2 _36514_ (.A(_08589_),
    .B(_08591_),
    .Y(_08592_));
 sky130_fd_sc_hd__a21oi_2 _36515_ (.A1(_08396_),
    .A2(_08405_),
    .B1(_08402_),
    .Y(_08593_));
 sky130_fd_sc_hd__or2_2 _36516_ (.A(_08592_),
    .B(_08593_),
    .X(_08594_));
 sky130_fd_sc_hd__nand2_2 _36517_ (.A(_08592_),
    .B(_08593_),
    .Y(_08595_));
 sky130_fd_sc_hd__nand2_2 _36518_ (.A(_08594_),
    .B(_08595_),
    .Y(_08596_));
 sky130_fd_sc_hd__o21a_2 _36519_ (.A1(_08395_),
    .A2(_08406_),
    .B1(_08408_),
    .X(_08597_));
 sky130_fd_sc_hd__nor2_2 _36520_ (.A(_08596_),
    .B(_08597_),
    .Y(_08598_));
 sky130_fd_sc_hd__and2_2 _36521_ (.A(_08596_),
    .B(_08597_),
    .X(_08599_));
 sky130_fd_sc_hd__or2_2 _36522_ (.A(_08598_),
    .B(_08599_),
    .X(_08600_));
 sky130_fd_sc_hd__a21oi_2 _36523_ (.A1(_08419_),
    .A2(_08420_),
    .B1(_08417_),
    .Y(_08602_));
 sky130_fd_sc_hd__and3_2 _36524_ (.A(_06413_),
    .B(_04781_),
    .C(_08416_),
    .X(_08603_));
 sky130_fd_sc_hd__a21oi_2 _36525_ (.A1(_06413_),
    .A2(_04781_),
    .B1(_08416_),
    .Y(_08604_));
 sky130_fd_sc_hd__nor2_2 _36526_ (.A(_08603_),
    .B(_08604_),
    .Y(_08605_));
 sky130_fd_sc_hd__nor2_2 _36527_ (.A(_05979_),
    .B(_05440_),
    .Y(_08606_));
 sky130_fd_sc_hd__xor2_2 _36528_ (.A(_08605_),
    .B(_08606_),
    .X(_08607_));
 sky130_fd_sc_hd__nand2_2 _36529_ (.A(_06983_),
    .B(_00567_),
    .Y(_08608_));
 sky130_fd_sc_hd__nand2_2 _36530_ (.A(_05450_),
    .B(_06983_),
    .Y(_08609_));
 sky130_fd_sc_hd__o21a_2 _36531_ (.A1(_06816_),
    .A2(_02311_),
    .B1(_08609_),
    .X(_08610_));
 sky130_fd_sc_hd__o21bai_2 _36532_ (.A1(_08422_),
    .A2(_08608_),
    .B1_N(_08610_),
    .Y(_08611_));
 sky130_fd_sc_hd__buf_1 _36533_ (.A(_03327_),
    .X(_08613_));
 sky130_fd_sc_hd__nand2_2 _36534_ (.A(_04138_),
    .B(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__xnor2_2 _36535_ (.A(_08611_),
    .B(_08614_),
    .Y(_08615_));
 sky130_fd_sc_hd__o21a_2 _36536_ (.A1(_08188_),
    .A2(_08422_),
    .B1(_08424_),
    .X(_08616_));
 sky130_fd_sc_hd__xor2_2 _36537_ (.A(_08615_),
    .B(_08616_),
    .X(_08617_));
 sky130_fd_sc_hd__nand2_2 _36538_ (.A(_08607_),
    .B(_08617_),
    .Y(_08618_));
 sky130_fd_sc_hd__or2_2 _36539_ (.A(_08607_),
    .B(_08617_),
    .X(_08619_));
 sky130_fd_sc_hd__nand2_2 _36540_ (.A(_08618_),
    .B(_08619_),
    .Y(_08620_));
 sky130_fd_sc_hd__a21oi_2 _36541_ (.A1(_08429_),
    .A2(_08432_),
    .B1(_08620_),
    .Y(_08621_));
 sky130_fd_sc_hd__and3_2 _36542_ (.A(_08429_),
    .B(_08432_),
    .C(_08620_),
    .X(_08622_));
 sky130_fd_sc_hd__nor2_2 _36543_ (.A(_08621_),
    .B(_08622_),
    .Y(_08624_));
 sky130_fd_sc_hd__xnor2_2 _36544_ (.A(_08602_),
    .B(_08624_),
    .Y(_08625_));
 sky130_fd_sc_hd__inv_2 _36545_ (.A(_08625_),
    .Y(_08626_));
 sky130_fd_sc_hd__or2_2 _36546_ (.A(_08600_),
    .B(_08626_),
    .X(_08627_));
 sky130_fd_sc_hd__nand2_2 _36547_ (.A(_08600_),
    .B(_08626_),
    .Y(_08628_));
 sky130_fd_sc_hd__o21ai_2 _36548_ (.A1(_08413_),
    .A2(_08439_),
    .B1(_08411_),
    .Y(_08629_));
 sky130_fd_sc_hd__and3_2 _36549_ (.A(_08627_),
    .B(_08628_),
    .C(_08629_),
    .X(_08630_));
 sky130_fd_sc_hd__a21oi_2 _36550_ (.A1(_08627_),
    .A2(_08628_),
    .B1(_08629_),
    .Y(_08631_));
 sky130_fd_sc_hd__nor2_2 _36551_ (.A(_08630_),
    .B(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__xnor2_2 _36552_ (.A(_08576_),
    .B(_08632_),
    .Y(_08633_));
 sky130_fd_sc_hd__a21boi_2 _36553_ (.A1(_08390_),
    .A2(_08443_),
    .B1_N(_08389_),
    .Y(_08635_));
 sky130_fd_sc_hd__xnor2_2 _36554_ (.A(_08633_),
    .B(_08635_),
    .Y(_08636_));
 sky130_fd_sc_hd__a21oi_2 _36555_ (.A1(_08414_),
    .A2(_08438_),
    .B1(_08435_),
    .Y(_08637_));
 sky130_fd_sc_hd__xnor2_2 _36556_ (.A(_08441_),
    .B(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__xor2_2 _36557_ (.A(_08636_),
    .B(_08638_),
    .X(_08639_));
 sky130_fd_sc_hd__a21boi_2 _36558_ (.A1(_08447_),
    .A2(_08453_),
    .B1_N(_08446_),
    .Y(_08640_));
 sky130_fd_sc_hd__nor2_2 _36559_ (.A(_08639_),
    .B(_08640_),
    .Y(_08641_));
 sky130_fd_sc_hd__and2_2 _36560_ (.A(_08639_),
    .B(_08640_),
    .X(_08642_));
 sky130_fd_sc_hd__nor2_2 _36561_ (.A(_08641_),
    .B(_08642_),
    .Y(_08643_));
 sky130_fd_sc_hd__xnor2_2 _36562_ (.A(_08560_),
    .B(_08643_),
    .Y(_08644_));
 sky130_fd_sc_hd__inv_2 _36563_ (.A(_08456_),
    .Y(_08646_));
 sky130_fd_sc_hd__nor2_2 _36564_ (.A(_08646_),
    .B(_08458_),
    .Y(_08647_));
 sky130_fd_sc_hd__xnor2_2 _36565_ (.A(_08644_),
    .B(_08647_),
    .Y(_08648_));
 sky130_fd_sc_hd__or4_2 _36566_ (.A(_08050_),
    .B(_08252_),
    .C(_08461_),
    .D(_08462_),
    .X(_08649_));
 sky130_fd_sc_hd__a211o_2 _36567_ (.A1(_07691_),
    .A2(_07694_),
    .B1(_08649_),
    .C1(_07807_),
    .X(_08650_));
 sky130_fd_sc_hd__and3_2 _36568_ (.A(_07796_),
    .B(_07799_),
    .C(_08048_),
    .X(_08651_));
 sky130_fd_sc_hd__a21o_2 _36569_ (.A1(_07805_),
    .A2(_08159_),
    .B1(_08651_),
    .X(_08652_));
 sky130_fd_sc_hd__or2_2 _36570_ (.A(_08366_),
    .B(_08462_),
    .X(_08653_));
 sky130_fd_sc_hd__inv_2 _36571_ (.A(_08461_),
    .Y(_08654_));
 sky130_fd_sc_hd__o311a_2 _36572_ (.A1(_08252_),
    .A2(_08462_),
    .A3(_08652_),
    .B1(_08653_),
    .C1(_08654_),
    .X(_08655_));
 sky130_fd_sc_hd__and2_2 _36573_ (.A(_08650_),
    .B(_08655_),
    .X(_08657_));
 sky130_fd_sc_hd__xnor2_2 _36574_ (.A(_08648_),
    .B(_08657_),
    .Y(_08658_));
 sky130_fd_sc_hd__and3_2 _36575_ (.A(iY[53]),
    .B(iX[63]),
    .C(_08468_),
    .X(_08659_));
 sky130_fd_sc_hd__a21o_2 _36576_ (.A1(iY[53]),
    .A2(iX[63]),
    .B1(_08468_),
    .X(_08660_));
 sky130_fd_sc_hd__and2b_2 _36577_ (.A_N(_08659_),
    .B(_08660_),
    .X(_08661_));
 sky130_fd_sc_hd__nand2_2 _36578_ (.A(iY[55]),
    .B(iX[61]),
    .Y(_08662_));
 sky130_fd_sc_hd__xnor2_2 _36579_ (.A(_08661_),
    .B(_08662_),
    .Y(_08663_));
 sky130_fd_sc_hd__inv_2 _36580_ (.A(_08663_),
    .Y(_08664_));
 sky130_fd_sc_hd__inv_2 _36581_ (.A(_08516_),
    .Y(_08665_));
 sky130_fd_sc_hd__and2b_2 _36582_ (.A_N(_08498_),
    .B(_08504_),
    .X(_08666_));
 sky130_fd_sc_hd__a21oi_2 _36583_ (.A1(_08467_),
    .A2(_08475_),
    .B1(_08255_),
    .Y(_08668_));
 sky130_fd_sc_hd__o21ba_2 _36584_ (.A1(_08500_),
    .A2(_08502_),
    .B1_N(_08499_),
    .X(_08669_));
 sky130_fd_sc_hd__and4_2 _36585_ (.A(iY[56]),
    .B(iY[57]),
    .C(iX[59]),
    .D(iX[60]),
    .X(_08670_));
 sky130_fd_sc_hd__a22oi_2 _36586_ (.A1(iY[57]),
    .A2(iX[59]),
    .B1(iX[60]),
    .B2(iY[56]),
    .Y(_08671_));
 sky130_fd_sc_hd__nor2_2 _36587_ (.A(_08670_),
    .B(_08671_),
    .Y(_08672_));
 sky130_fd_sc_hd__a21oi_2 _36588_ (.A1(iX[58]),
    .A2(iY[58]),
    .B1(_08672_),
    .Y(_08673_));
 sky130_fd_sc_hd__and3_2 _36589_ (.A(iX[58]),
    .B(iY[58]),
    .C(_08672_),
    .X(_08674_));
 sky130_fd_sc_hd__nor2_2 _36590_ (.A(_08673_),
    .B(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__o21a_2 _36591_ (.A1(_08469_),
    .A2(_08474_),
    .B1(_08675_),
    .X(_08676_));
 sky130_fd_sc_hd__nor3_2 _36592_ (.A(_08469_),
    .B(_08474_),
    .C(_08675_),
    .Y(_08677_));
 sky130_fd_sc_hd__nor2_2 _36593_ (.A(_08676_),
    .B(_08677_),
    .Y(_08679_));
 sky130_fd_sc_hd__xnor2_2 _36594_ (.A(_08669_),
    .B(_08679_),
    .Y(_08680_));
 sky130_fd_sc_hd__xnor2_2 _36595_ (.A(_08668_),
    .B(_08680_),
    .Y(_08681_));
 sky130_fd_sc_hd__o21ai_2 _36596_ (.A1(_08666_),
    .A2(_08506_),
    .B1(_08681_),
    .Y(_08682_));
 sky130_fd_sc_hd__or3_2 _36597_ (.A(_08666_),
    .B(_08506_),
    .C(_08681_),
    .X(_08683_));
 sky130_fd_sc_hd__or2b_2 _36598_ (.A(_08509_),
    .B_N(_08511_),
    .X(_08684_));
 sky130_fd_sc_hd__and3_2 _36599_ (.A(_08682_),
    .B(_08683_),
    .C(_08684_),
    .X(_08685_));
 sky130_fd_sc_hd__inv_2 _36600_ (.A(_08685_),
    .Y(_08686_));
 sky130_fd_sc_hd__a21o_2 _36601_ (.A1(_08682_),
    .A2(_08683_),
    .B1(_08684_),
    .X(_08687_));
 sky130_fd_sc_hd__or2b_2 _36602_ (.A(_08484_),
    .B_N(_08483_),
    .X(_08688_));
 sky130_fd_sc_hd__and4_2 _36603_ (.A(iX[56]),
    .B(iX[57]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_08690_));
 sky130_fd_sc_hd__a22oi_2 _36604_ (.A1(iX[57]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[56]),
    .Y(_08691_));
 sky130_fd_sc_hd__nor2_2 _36605_ (.A(_08690_),
    .B(_08691_),
    .Y(_08692_));
 sky130_fd_sc_hd__nand2_2 _36606_ (.A(iX[55]),
    .B(iY[61]),
    .Y(_08693_));
 sky130_fd_sc_hd__xnor2_2 _36607_ (.A(_08692_),
    .B(_08693_),
    .Y(_08694_));
 sky130_fd_sc_hd__o21ba_2 _36608_ (.A1(_08479_),
    .A2(_08482_),
    .B1_N(_08478_),
    .X(_08695_));
 sky130_fd_sc_hd__xnor2_2 _36609_ (.A(_08694_),
    .B(_08695_),
    .Y(_08696_));
 sky130_fd_sc_hd__and2_2 _36610_ (.A(iX[54]),
    .B(iY[62]),
    .X(_08697_));
 sky130_fd_sc_hd__or2_2 _36611_ (.A(_08696_),
    .B(_08697_),
    .X(_08698_));
 sky130_fd_sc_hd__nand2_2 _36612_ (.A(_08696_),
    .B(_08697_),
    .Y(_08699_));
 sky130_fd_sc_hd__nand2_2 _36613_ (.A(_08698_),
    .B(_08699_),
    .Y(_08701_));
 sky130_fd_sc_hd__a21oi_2 _36614_ (.A1(_08688_),
    .A2(_08488_),
    .B1(_08701_),
    .Y(_08702_));
 sky130_fd_sc_hd__and3_2 _36615_ (.A(_08688_),
    .B(_08488_),
    .C(_08701_),
    .X(_08703_));
 sky130_fd_sc_hd__nor2_2 _36616_ (.A(_08702_),
    .B(_08703_),
    .Y(_08704_));
 sky130_fd_sc_hd__nand2_2 _36617_ (.A(iX[53]),
    .B(iY[63]),
    .Y(_08705_));
 sky130_fd_sc_hd__xnor2_2 _36618_ (.A(_08704_),
    .B(_08705_),
    .Y(_08706_));
 sky130_fd_sc_hd__a21oi_2 _36619_ (.A1(_08686_),
    .A2(_08687_),
    .B1(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__and3_2 _36620_ (.A(_08686_),
    .B(_08687_),
    .C(_08706_),
    .X(_08708_));
 sky130_fd_sc_hd__a211o_2 _36621_ (.A1(_08513_),
    .A2(_08665_),
    .B1(_08707_),
    .C1(_08708_),
    .X(_08709_));
 sky130_fd_sc_hd__o211ai_2 _36622_ (.A1(_08707_),
    .A2(_08708_),
    .B1(_08513_),
    .C1(_08665_),
    .Y(_08710_));
 sky130_fd_sc_hd__nand2_2 _36623_ (.A(_08709_),
    .B(_08710_),
    .Y(_08712_));
 sky130_fd_sc_hd__nor2_2 _36624_ (.A(_08664_),
    .B(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__and2_2 _36625_ (.A(_08664_),
    .B(_08712_),
    .X(_08714_));
 sky130_fd_sc_hd__or2_2 _36626_ (.A(_08713_),
    .B(_08714_),
    .X(_08715_));
 sky130_fd_sc_hd__or2_2 _36627_ (.A(_08522_),
    .B(_08715_),
    .X(_08716_));
 sky130_fd_sc_hd__nand2_2 _36628_ (.A(_08522_),
    .B(_08715_),
    .Y(_08717_));
 sky130_fd_sc_hd__and2_2 _36629_ (.A(_08716_),
    .B(_08717_),
    .X(_08718_));
 sky130_fd_sc_hd__o21ai_2 _36630_ (.A1(_08518_),
    .A2(_08520_),
    .B1(_08718_),
    .Y(_08719_));
 sky130_fd_sc_hd__or3_2 _36631_ (.A(_08518_),
    .B(_08520_),
    .C(_08718_),
    .X(_08720_));
 sky130_fd_sc_hd__and2_2 _36632_ (.A(_08719_),
    .B(_08720_),
    .X(_08721_));
 sky130_fd_sc_hd__o21ai_2 _36633_ (.A1(_08524_),
    .A2(_08528_),
    .B1(_08721_),
    .Y(_08723_));
 sky130_fd_sc_hd__or3_2 _36634_ (.A(_08524_),
    .B(_08528_),
    .C(_08721_),
    .X(_08724_));
 sky130_fd_sc_hd__nand2_2 _36635_ (.A(_08723_),
    .B(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__a31o_2 _36636_ (.A1(iX[52]),
    .A2(iY[63]),
    .A3(_08493_),
    .B1(_08490_),
    .X(_08726_));
 sky130_fd_sc_hd__xnor2_2 _36637_ (.A(_08725_),
    .B(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__o21ai_2 _36638_ (.A1(_08530_),
    .A2(_08532_),
    .B1(_08727_),
    .Y(_08728_));
 sky130_fd_sc_hd__or3_2 _36639_ (.A(_08530_),
    .B(_08532_),
    .C(_08727_),
    .X(_08729_));
 sky130_fd_sc_hd__nand2_2 _36640_ (.A(_08728_),
    .B(_08729_),
    .Y(_08730_));
 sky130_fd_sc_hd__nand2_2 _36641_ (.A(_08340_),
    .B(_08538_),
    .Y(_08731_));
 sky130_fd_sc_hd__a2111o_2 _36642_ (.A1(_07907_),
    .A2(_07909_),
    .B1(_08144_),
    .C1(_08731_),
    .D1(_07905_),
    .X(_08732_));
 sky130_fd_sc_hd__nand2_2 _36643_ (.A(_08337_),
    .B(_08535_),
    .Y(_08734_));
 sky130_fd_sc_hd__o211a_2 _36644_ (.A1(_08341_),
    .A2(_08731_),
    .B1(_08734_),
    .C1(_08537_),
    .X(_08735_));
 sky130_fd_sc_hd__and2_2 _36645_ (.A(_08732_),
    .B(_08735_),
    .X(_08736_));
 sky130_fd_sc_hd__xnor2_2 _36646_ (.A(_08730_),
    .B(_08736_),
    .Y(_08737_));
 sky130_fd_sc_hd__xnor2_2 _36647_ (.A(_08658_),
    .B(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__and2_2 _36648_ (.A(_16890_),
    .B(_08738_),
    .X(_08739_));
 sky130_fd_sc_hd__nor2_2 _36649_ (.A(_16890_),
    .B(_08738_),
    .Y(_08740_));
 sky130_fd_sc_hd__or2_2 _36650_ (.A(_08739_),
    .B(_08740_),
    .X(_08741_));
 sky130_fd_sc_hd__a21boi_2 _36651_ (.A1(_16809_),
    .A2(_08541_),
    .B1_N(_08542_),
    .Y(_08742_));
 sky130_fd_sc_hd__nor2_2 _36652_ (.A(_08741_),
    .B(_08742_),
    .Y(_08743_));
 sky130_fd_sc_hd__and2_2 _36653_ (.A(_08741_),
    .B(_08742_),
    .X(_08745_));
 sky130_fd_sc_hd__nor2_2 _36654_ (.A(_08743_),
    .B(_08745_),
    .Y(_08746_));
 sky130_fd_sc_hd__o311a_2 _36655_ (.A1(_08347_),
    .A2(_08349_),
    .A3(_08546_),
    .B1(_08548_),
    .C1(_08358_),
    .X(_08747_));
 sky130_fd_sc_hd__a21o_2 _36656_ (.A1(_08352_),
    .A2(_08548_),
    .B1(_08546_),
    .X(_08748_));
 sky130_fd_sc_hd__a21oi_4 _36657_ (.A1(_08355_),
    .A2(_08747_),
    .B1(_08748_),
    .Y(_08749_));
 sky130_fd_sc_hd__xor2_2 _36658_ (.A(_08746_),
    .B(_08749_),
    .X(_08750_));
 sky130_fd_sc_hd__nand2_2 _36659_ (.A(_17171_),
    .B(_08750_),
    .Y(_08751_));
 sky130_fd_sc_hd__or2_2 _36660_ (.A(_17171_),
    .B(_08750_),
    .X(_08752_));
 sky130_fd_sc_hd__and2_2 _36661_ (.A(_08751_),
    .B(_08752_),
    .X(_08753_));
 sky130_fd_sc_hd__and2b_2 _36662_ (.A_N(_08559_),
    .B(_08753_),
    .X(_08754_));
 sky130_fd_sc_hd__and2b_2 _36663_ (.A_N(_08753_),
    .B(_08559_),
    .X(_08756_));
 sky130_fd_sc_hd__nor2_2 _36664_ (.A(_08754_),
    .B(_08756_),
    .Y(oO[84]));
 sky130_fd_sc_hd__and2b_2 _36665_ (.A_N(_08658_),
    .B(_08737_),
    .X(_08757_));
 sky130_fd_sc_hd__nand2_2 _36666_ (.A(_08225_),
    .B(_08227_),
    .Y(_08758_));
 sky130_fd_sc_hd__or3b_2 _36667_ (.A(_08637_),
    .B(_08440_),
    .C_N(_08758_),
    .X(_08759_));
 sky130_fd_sc_hd__nor2_2 _36668_ (.A(_08570_),
    .B(_08574_),
    .Y(_08760_));
 sky130_fd_sc_hd__nand2_2 _36669_ (.A(_06813_),
    .B(_06783_),
    .Y(_08761_));
 sky130_fd_sc_hd__a21bo_2 _36670_ (.A1(_08562_),
    .A2(_08569_),
    .B1_N(_08561_),
    .X(_08762_));
 sky130_fd_sc_hd__buf_1 _36671_ (.A(_05533_),
    .X(_08763_));
 sky130_fd_sc_hd__o22a_2 _36672_ (.A1(_05979_),
    .A2(_06786_),
    .B1(_08164_),
    .B2(_05978_),
    .X(_08764_));
 sky130_fd_sc_hd__a31o_2 _36673_ (.A1(_06411_),
    .A2(_05507_),
    .A3(_08763_),
    .B1(_08764_),
    .X(_08766_));
 sky130_fd_sc_hd__xnor2_2 _36674_ (.A(_08762_),
    .B(_08766_),
    .Y(_08767_));
 sky130_fd_sc_hd__xnor2_2 _36675_ (.A(_08761_),
    .B(_08767_),
    .Y(_08768_));
 sky130_fd_sc_hd__xnor2_2 _36676_ (.A(_08760_),
    .B(_08768_),
    .Y(_08769_));
 sky130_fd_sc_hd__nor2_2 _36677_ (.A(_08600_),
    .B(_08626_),
    .Y(_08770_));
 sky130_fd_sc_hd__or3_2 _36678_ (.A(_08580_),
    .B(_08585_),
    .C(_08586_),
    .X(_08771_));
 sky130_fd_sc_hd__nor2_2 _36679_ (.A(_18344_),
    .B(_06797_),
    .Y(_08772_));
 sky130_fd_sc_hd__and3_2 _36680_ (.A(_07039_),
    .B(_03994_),
    .C(_08772_),
    .X(_08773_));
 sky130_fd_sc_hd__o22a_2 _36681_ (.A1(_18344_),
    .A2(_08582_),
    .B1(_06797_),
    .B2(_06491_),
    .X(_08774_));
 sky130_fd_sc_hd__nor2_2 _36682_ (.A(_08773_),
    .B(_08774_),
    .Y(_08775_));
 sky130_fd_sc_hd__and3_2 _36683_ (.A(_06484_),
    .B(_07472_),
    .C(_08775_),
    .X(_08777_));
 sky130_fd_sc_hd__a21oi_2 _36684_ (.A1(_06484_),
    .A2(_07472_),
    .B1(_08775_),
    .Y(_08778_));
 sky130_fd_sc_hd__or2_2 _36685_ (.A(_08777_),
    .B(_08778_),
    .X(_08779_));
 sky130_fd_sc_hd__xnor2_2 _36686_ (.A(_08573_),
    .B(_08779_),
    .Y(_08780_));
 sky130_fd_sc_hd__o21ai_2 _36687_ (.A1(_08581_),
    .A2(_08585_),
    .B1(_08780_),
    .Y(_08781_));
 sky130_fd_sc_hd__or3_2 _36688_ (.A(_08581_),
    .B(_08585_),
    .C(_08780_),
    .X(_08782_));
 sky130_fd_sc_hd__nand2_2 _36689_ (.A(_08781_),
    .B(_08782_),
    .Y(_08783_));
 sky130_fd_sc_hd__a21oi_2 _36690_ (.A1(_08771_),
    .A2(_08589_),
    .B1(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__and3_2 _36691_ (.A(_08771_),
    .B(_08589_),
    .C(_08783_),
    .X(_08785_));
 sky130_fd_sc_hd__or2_2 _36692_ (.A(_08784_),
    .B(_08785_),
    .X(_08786_));
 sky130_fd_sc_hd__nor2_2 _36693_ (.A(_08594_),
    .B(_08786_),
    .Y(_08788_));
 sky130_fd_sc_hd__and2_2 _36694_ (.A(_08594_),
    .B(_08786_),
    .X(_08789_));
 sky130_fd_sc_hd__or2_2 _36695_ (.A(_08788_),
    .B(_08789_),
    .X(_08790_));
 sky130_fd_sc_hd__a21oi_2 _36696_ (.A1(_08605_),
    .A2(_08606_),
    .B1(_08603_),
    .Y(_08791_));
 sky130_fd_sc_hd__or2_2 _36697_ (.A(_08615_),
    .B(_08616_),
    .X(_08792_));
 sky130_fd_sc_hd__nor2_2 _36698_ (.A(_05522_),
    .B(_07252_),
    .Y(_08793_));
 sky130_fd_sc_hd__and3_2 _36699_ (.A(_06413_),
    .B(_07007_),
    .C(_08793_),
    .X(_08794_));
 sky130_fd_sc_hd__buf_1 _36700_ (.A(_07252_),
    .X(_08795_));
 sky130_fd_sc_hd__o22a_2 _36701_ (.A1(_05522_),
    .A2(_04782_),
    .B1(_08795_),
    .B2(_05504_),
    .X(_08796_));
 sky130_fd_sc_hd__nor2_2 _36702_ (.A(_08794_),
    .B(_08796_),
    .Y(_08797_));
 sky130_fd_sc_hd__nor2_2 _36703_ (.A(_04862_),
    .B(_05441_),
    .Y(_08799_));
 sky130_fd_sc_hd__xor2_2 _36704_ (.A(_08797_),
    .B(_08799_),
    .X(_08800_));
 sky130_fd_sc_hd__nand2_2 _36705_ (.A(_05450_),
    .B(_07461_),
    .Y(_08801_));
 sky130_fd_sc_hd__xnor2_2 _36706_ (.A(_08608_),
    .B(_08801_),
    .Y(_08802_));
 sky130_fd_sc_hd__nand2_2 _36707_ (.A(_06822_),
    .B(_08613_),
    .Y(_08803_));
 sky130_fd_sc_hd__xnor2_2 _36708_ (.A(_08802_),
    .B(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__o22a_2 _36709_ (.A1(_08422_),
    .A2(_08608_),
    .B1(_08610_),
    .B2(_08614_),
    .X(_08805_));
 sky130_fd_sc_hd__or2_2 _36710_ (.A(_08804_),
    .B(_08805_),
    .X(_08806_));
 sky130_fd_sc_hd__nand2_2 _36711_ (.A(_08804_),
    .B(_08805_),
    .Y(_08807_));
 sky130_fd_sc_hd__and2_2 _36712_ (.A(_08806_),
    .B(_08807_),
    .X(_08808_));
 sky130_fd_sc_hd__nand2_2 _36713_ (.A(_08800_),
    .B(_08808_),
    .Y(_08810_));
 sky130_fd_sc_hd__or2_2 _36714_ (.A(_08800_),
    .B(_08808_),
    .X(_08811_));
 sky130_fd_sc_hd__nand2_2 _36715_ (.A(_08810_),
    .B(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__a21oi_2 _36716_ (.A1(_08792_),
    .A2(_08618_),
    .B1(_08812_),
    .Y(_08813_));
 sky130_fd_sc_hd__and3_2 _36717_ (.A(_08792_),
    .B(_08618_),
    .C(_08812_),
    .X(_08814_));
 sky130_fd_sc_hd__nor2_2 _36718_ (.A(_08813_),
    .B(_08814_),
    .Y(_08815_));
 sky130_fd_sc_hd__xnor2_2 _36719_ (.A(_08791_),
    .B(_08815_),
    .Y(_08816_));
 sky130_fd_sc_hd__xnor2_2 _36720_ (.A(_08790_),
    .B(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__o21a_2 _36721_ (.A1(_08598_),
    .A2(_08770_),
    .B1(_08817_),
    .X(_08818_));
 sky130_fd_sc_hd__nor3_2 _36722_ (.A(_08598_),
    .B(_08770_),
    .C(_08817_),
    .Y(_08819_));
 sky130_fd_sc_hd__nor2_2 _36723_ (.A(_08818_),
    .B(_08819_),
    .Y(_08821_));
 sky130_fd_sc_hd__xnor2_2 _36724_ (.A(_08769_),
    .B(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__and3_2 _36725_ (.A(_08380_),
    .B(_08385_),
    .C(_08386_),
    .X(_08823_));
 sky130_fd_sc_hd__and2_2 _36726_ (.A(_08576_),
    .B(_08632_),
    .X(_08824_));
 sky130_fd_sc_hd__a21oi_2 _36727_ (.A1(_08823_),
    .A2(_08575_),
    .B1(_08824_),
    .Y(_08825_));
 sky130_fd_sc_hd__xnor2_2 _36728_ (.A(_08822_),
    .B(_08825_),
    .Y(_08826_));
 sky130_fd_sc_hd__and2b_2 _36729_ (.A_N(_08602_),
    .B(_08624_),
    .X(_08827_));
 sky130_fd_sc_hd__o21ai_2 _36730_ (.A1(_08621_),
    .A2(_08827_),
    .B1(_08630_),
    .Y(_08828_));
 sky130_fd_sc_hd__or3_2 _36731_ (.A(_08621_),
    .B(_08827_),
    .C(_08630_),
    .X(_08829_));
 sky130_fd_sc_hd__and2_2 _36732_ (.A(_08828_),
    .B(_08829_),
    .X(_08830_));
 sky130_fd_sc_hd__xnor2_2 _36733_ (.A(_08826_),
    .B(_08830_),
    .Y(_08832_));
 sky130_fd_sc_hd__or2b_2 _36734_ (.A(_08636_),
    .B_N(_08638_),
    .X(_08833_));
 sky130_fd_sc_hd__o21ai_2 _36735_ (.A1(_08633_),
    .A2(_08635_),
    .B1(_08833_),
    .Y(_08834_));
 sky130_fd_sc_hd__xor2_2 _36736_ (.A(_08832_),
    .B(_08834_),
    .X(_08835_));
 sky130_fd_sc_hd__xnor2_2 _36737_ (.A(_08759_),
    .B(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__a21oi_2 _36738_ (.A1(_08560_),
    .A2(_08643_),
    .B1(_08641_),
    .Y(_08837_));
 sky130_fd_sc_hd__xor2_2 _36739_ (.A(_08836_),
    .B(_08837_),
    .X(_08838_));
 sky130_fd_sc_hd__nor2_2 _36740_ (.A(_08644_),
    .B(_08647_),
    .Y(_08839_));
 sky130_fd_sc_hd__o21ba_2 _36741_ (.A1(_08648_),
    .A2(_08657_),
    .B1_N(_08839_),
    .X(_08840_));
 sky130_fd_sc_hd__xnor2_2 _36742_ (.A(_08838_),
    .B(_08840_),
    .Y(_08841_));
 sky130_fd_sc_hd__or2b_2 _36743_ (.A(_08725_),
    .B_N(_08726_),
    .X(_08843_));
 sky130_fd_sc_hd__a22oi_2 _36744_ (.A1(iY[55]),
    .A2(iX[62]),
    .B1(iX[63]),
    .B2(iY[54]),
    .Y(_08844_));
 sky130_fd_sc_hd__and3_2 _36745_ (.A(iY[55]),
    .B(iX[63]),
    .C(_08468_),
    .X(_08845_));
 sky130_fd_sc_hd__or2_2 _36746_ (.A(_08844_),
    .B(_08845_),
    .X(_08846_));
 sky130_fd_sc_hd__a31o_2 _36747_ (.A1(iY[55]),
    .A2(iX[61]),
    .A3(_08660_),
    .B1(_08659_),
    .X(_08847_));
 sky130_fd_sc_hd__nand4_2 _36748_ (.A(iY[56]),
    .B(iY[57]),
    .C(iX[60]),
    .D(iX[61]),
    .Y(_08848_));
 sky130_fd_sc_hd__a22o_2 _36749_ (.A1(iY[57]),
    .A2(iX[60]),
    .B1(iX[61]),
    .B2(iY[56]),
    .X(_08849_));
 sky130_fd_sc_hd__nand2_2 _36750_ (.A(_08848_),
    .B(_08849_),
    .Y(_08850_));
 sky130_fd_sc_hd__nand2_2 _36751_ (.A(iY[58]),
    .B(iX[59]),
    .Y(_08851_));
 sky130_fd_sc_hd__xor2_2 _36752_ (.A(_08850_),
    .B(_08851_),
    .X(_08852_));
 sky130_fd_sc_hd__xor2_2 _36753_ (.A(_08847_),
    .B(_08852_),
    .X(_08854_));
 sky130_fd_sc_hd__or3_2 _36754_ (.A(_08670_),
    .B(_08674_),
    .C(_08854_),
    .X(_08855_));
 sky130_fd_sc_hd__o21ai_2 _36755_ (.A1(_08670_),
    .A2(_08674_),
    .B1(_08854_),
    .Y(_08856_));
 sky130_fd_sc_hd__nand2_2 _36756_ (.A(_08855_),
    .B(_08856_),
    .Y(_08857_));
 sky130_fd_sc_hd__o21ba_2 _36757_ (.A1(_08669_),
    .A2(_08677_),
    .B1_N(_08676_),
    .X(_08858_));
 sky130_fd_sc_hd__or2_2 _36758_ (.A(_08857_),
    .B(_08858_),
    .X(_08859_));
 sky130_fd_sc_hd__nand2_2 _36759_ (.A(_08857_),
    .B(_08858_),
    .Y(_08860_));
 sky130_fd_sc_hd__nand2_2 _36760_ (.A(_08859_),
    .B(_08860_),
    .Y(_08861_));
 sky130_fd_sc_hd__inv_2 _36761_ (.A(_08680_),
    .Y(_08862_));
 sky130_fd_sc_hd__o21a_2 _36762_ (.A1(_08668_),
    .A2(_08862_),
    .B1(_08682_),
    .X(_08863_));
 sky130_fd_sc_hd__nor2_2 _36763_ (.A(_08861_),
    .B(_08863_),
    .Y(_08865_));
 sky130_fd_sc_hd__and2_2 _36764_ (.A(_08861_),
    .B(_08863_),
    .X(_08866_));
 sky130_fd_sc_hd__nor2_2 _36765_ (.A(_08865_),
    .B(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__or2b_2 _36766_ (.A(_08695_),
    .B_N(_08694_),
    .X(_08868_));
 sky130_fd_sc_hd__and4_2 _36767_ (.A(iX[57]),
    .B(iX[58]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_08869_));
 sky130_fd_sc_hd__a22oi_2 _36768_ (.A1(iX[58]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[57]),
    .Y(_08870_));
 sky130_fd_sc_hd__nor2_2 _36769_ (.A(_08869_),
    .B(_08870_),
    .Y(_08871_));
 sky130_fd_sc_hd__nand2_2 _36770_ (.A(iX[56]),
    .B(iY[61]),
    .Y(_08872_));
 sky130_fd_sc_hd__xnor2_2 _36771_ (.A(_08871_),
    .B(_08872_),
    .Y(_08873_));
 sky130_fd_sc_hd__o21ba_2 _36772_ (.A1(_08691_),
    .A2(_08693_),
    .B1_N(_08690_),
    .X(_08874_));
 sky130_fd_sc_hd__xnor2_2 _36773_ (.A(_08873_),
    .B(_08874_),
    .Y(_08876_));
 sky130_fd_sc_hd__and2_2 _36774_ (.A(iX[55]),
    .B(iY[62]),
    .X(_08877_));
 sky130_fd_sc_hd__or2_2 _36775_ (.A(_08876_),
    .B(_08877_),
    .X(_08878_));
 sky130_fd_sc_hd__nand2_2 _36776_ (.A(_08876_),
    .B(_08877_),
    .Y(_08879_));
 sky130_fd_sc_hd__nand2_2 _36777_ (.A(_08878_),
    .B(_08879_),
    .Y(_08880_));
 sky130_fd_sc_hd__a21oi_2 _36778_ (.A1(_08868_),
    .A2(_08699_),
    .B1(_08880_),
    .Y(_08881_));
 sky130_fd_sc_hd__and3_2 _36779_ (.A(_08868_),
    .B(_08699_),
    .C(_08880_),
    .X(_08882_));
 sky130_fd_sc_hd__nor2_2 _36780_ (.A(_08881_),
    .B(_08882_),
    .Y(_08883_));
 sky130_fd_sc_hd__nand2_2 _36781_ (.A(iX[54]),
    .B(iY[63]),
    .Y(_08884_));
 sky130_fd_sc_hd__xnor2_2 _36782_ (.A(_08883_),
    .B(_08884_),
    .Y(_08885_));
 sky130_fd_sc_hd__xor2_2 _36783_ (.A(_08867_),
    .B(_08885_),
    .X(_08887_));
 sky130_fd_sc_hd__o21a_2 _36784_ (.A1(_08685_),
    .A2(_08708_),
    .B1(_08887_),
    .X(_08888_));
 sky130_fd_sc_hd__nor2_2 _36785_ (.A(_08685_),
    .B(_08708_),
    .Y(_08889_));
 sky130_fd_sc_hd__and2b_2 _36786_ (.A_N(_08887_),
    .B(_08889_),
    .X(_08890_));
 sky130_fd_sc_hd__nor2_2 _36787_ (.A(_08888_),
    .B(_08890_),
    .Y(_08891_));
 sky130_fd_sc_hd__xnor2_2 _36788_ (.A(_08846_),
    .B(_08891_),
    .Y(_08892_));
 sky130_fd_sc_hd__or2_2 _36789_ (.A(_08713_),
    .B(_08892_),
    .X(_08893_));
 sky130_fd_sc_hd__nand2_2 _36790_ (.A(_08713_),
    .B(_08892_),
    .Y(_08894_));
 sky130_fd_sc_hd__nand2_2 _36791_ (.A(_08893_),
    .B(_08894_),
    .Y(_08895_));
 sky130_fd_sc_hd__xnor2_2 _36792_ (.A(_08709_),
    .B(_08895_),
    .Y(_08896_));
 sky130_fd_sc_hd__a21oi_2 _36793_ (.A1(_08716_),
    .A2(_08719_),
    .B1(_08896_),
    .Y(_08898_));
 sky130_fd_sc_hd__and3_2 _36794_ (.A(_08716_),
    .B(_08719_),
    .C(_08896_),
    .X(_08899_));
 sky130_fd_sc_hd__or2_2 _36795_ (.A(_08898_),
    .B(_08899_),
    .X(_08900_));
 sky130_fd_sc_hd__a31o_2 _36796_ (.A1(iX[53]),
    .A2(iY[63]),
    .A3(_08704_),
    .B1(_08702_),
    .X(_08901_));
 sky130_fd_sc_hd__xor2_2 _36797_ (.A(_08900_),
    .B(_08901_),
    .X(_08902_));
 sky130_fd_sc_hd__a21o_2 _36798_ (.A1(_08723_),
    .A2(_08843_),
    .B1(_08902_),
    .X(_08903_));
 sky130_fd_sc_hd__inv_2 _36799_ (.A(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__and3_2 _36800_ (.A(_08723_),
    .B(_08843_),
    .C(_08902_),
    .X(_08905_));
 sky130_fd_sc_hd__nor2_2 _36801_ (.A(_08904_),
    .B(_08905_),
    .Y(_08906_));
 sky130_fd_sc_hd__o21a_2 _36802_ (.A1(_08730_),
    .A2(_08736_),
    .B1(_08728_),
    .X(_08907_));
 sky130_fd_sc_hd__xnor2_2 _36803_ (.A(_08906_),
    .B(_08907_),
    .Y(_08909_));
 sky130_fd_sc_hd__xnor2_2 _36804_ (.A(_08841_),
    .B(_08909_),
    .Y(_08910_));
 sky130_fd_sc_hd__xor2_2 _36805_ (.A(_17259_),
    .B(_08910_),
    .X(_08911_));
 sky130_fd_sc_hd__o21a_2 _36806_ (.A1(_08757_),
    .A2(_08739_),
    .B1(_08911_),
    .X(_08912_));
 sky130_fd_sc_hd__or3_2 _36807_ (.A(_08757_),
    .B(_08739_),
    .C(_08911_),
    .X(_08913_));
 sky130_fd_sc_hd__and2b_2 _36808_ (.A_N(_08912_),
    .B(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__a21oi_2 _36809_ (.A1(_08746_),
    .A2(_08749_),
    .B1(_08743_),
    .Y(_08915_));
 sky130_fd_sc_hd__xnor2_2 _36810_ (.A(_08914_),
    .B(_08915_),
    .Y(_08916_));
 sky130_fd_sc_hd__and2_2 _36811_ (.A(_17376_),
    .B(_08916_),
    .X(_08917_));
 sky130_fd_sc_hd__nor2_2 _36812_ (.A(_17376_),
    .B(_08916_),
    .Y(_08918_));
 sky130_fd_sc_hd__nor2_2 _36813_ (.A(_08917_),
    .B(_08918_),
    .Y(_08920_));
 sky130_fd_sc_hd__a21oi_2 _36814_ (.A1(_17171_),
    .A2(_08750_),
    .B1(_08754_),
    .Y(_08921_));
 sky130_fd_sc_hd__xnor2_2 _36815_ (.A(_08920_),
    .B(_08921_),
    .Y(oO[85]));
 sky130_fd_sc_hd__and2b_2 _36816_ (.A_N(_08832_),
    .B(_08834_),
    .X(_08922_));
 sky130_fd_sc_hd__nor2_2 _36817_ (.A(_08759_),
    .B(_08835_),
    .Y(_08923_));
 sky130_fd_sc_hd__and3_2 _36818_ (.A(_06813_),
    .B(_06783_),
    .C(_08767_),
    .X(_08924_));
 sky130_fd_sc_hd__or2b_2 _36819_ (.A(_08563_),
    .B_N(_08569_),
    .X(_08925_));
 sky130_fd_sc_hd__buf_1 _36820_ (.A(_06399_),
    .X(_08926_));
 sky130_fd_sc_hd__or2_2 _36821_ (.A(_08926_),
    .B(_05976_),
    .X(_08927_));
 sky130_fd_sc_hd__a31o_2 _36822_ (.A1(_08561_),
    .A2(_08925_),
    .A3(_08927_),
    .B1(_08764_),
    .X(_08928_));
 sky130_fd_sc_hd__nor2_2 _36823_ (.A(_08926_),
    .B(_06814_),
    .Y(_08930_));
 sky130_fd_sc_hd__buf_1 _36824_ (.A(_06786_),
    .X(_08931_));
 sky130_fd_sc_hd__o22a_2 _36825_ (.A1(_04862_),
    .A2(_08931_),
    .B1(_08164_),
    .B2(_05500_),
    .X(_08932_));
 sky130_fd_sc_hd__nor2_2 _36826_ (.A(_08930_),
    .B(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__xnor2_2 _36827_ (.A(_08928_),
    .B(_08933_),
    .Y(_08934_));
 sky130_fd_sc_hd__xnor2_2 _36828_ (.A(_08924_),
    .B(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__and2b_2 _36829_ (.A_N(_08790_),
    .B(_08816_),
    .X(_08936_));
 sky130_fd_sc_hd__or3b_2 _36830_ (.A(_08777_),
    .B(_08778_),
    .C_N(_08573_),
    .X(_08937_));
 sky130_fd_sc_hd__and3_2 _36831_ (.A(_07039_),
    .B(_04905_),
    .C(_08772_),
    .X(_08938_));
 sky130_fd_sc_hd__a21oi_2 _36832_ (.A1(_07039_),
    .A2(_04905_),
    .B1(_08772_),
    .Y(_08939_));
 sky130_fd_sc_hd__nor2_2 _36833_ (.A(_08938_),
    .B(_08939_),
    .Y(_08941_));
 sky130_fd_sc_hd__and3_2 _36834_ (.A(_07279_),
    .B(_06154_),
    .C(_08941_),
    .X(_08942_));
 sky130_fd_sc_hd__a21oi_2 _36835_ (.A1(_07279_),
    .A2(_06154_),
    .B1(_08941_),
    .Y(_08943_));
 sky130_fd_sc_hd__nor2_2 _36836_ (.A(_08942_),
    .B(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__o21ai_2 _36837_ (.A1(_08773_),
    .A2(_08777_),
    .B1(_08944_),
    .Y(_08945_));
 sky130_fd_sc_hd__or3_2 _36838_ (.A(_08773_),
    .B(_08777_),
    .C(_08944_),
    .X(_08946_));
 sky130_fd_sc_hd__nand2_2 _36839_ (.A(_08945_),
    .B(_08946_),
    .Y(_08947_));
 sky130_fd_sc_hd__a21oi_2 _36840_ (.A1(_08937_),
    .A2(_08781_),
    .B1(_08947_),
    .Y(_08948_));
 sky130_fd_sc_hd__and3_2 _36841_ (.A(_08937_),
    .B(_08781_),
    .C(_08947_),
    .X(_08949_));
 sky130_fd_sc_hd__or3b_2 _36842_ (.A(_08948_),
    .B(_08949_),
    .C_N(_08784_),
    .X(_08950_));
 sky130_fd_sc_hd__or2_2 _36843_ (.A(_08948_),
    .B(_08949_),
    .X(_08952_));
 sky130_fd_sc_hd__or2b_2 _36844_ (.A(_08784_),
    .B_N(_08952_),
    .X(_08953_));
 sky130_fd_sc_hd__nand2_2 _36845_ (.A(_08950_),
    .B(_08953_),
    .Y(_08954_));
 sky130_fd_sc_hd__a21o_2 _36846_ (.A1(_08797_),
    .A2(_08799_),
    .B1(_08794_),
    .X(_08955_));
 sky130_fd_sc_hd__and3_2 _36847_ (.A(_06822_),
    .B(_04781_),
    .C(_08793_),
    .X(_08956_));
 sky130_fd_sc_hd__a21oi_2 _36848_ (.A1(_06822_),
    .A2(_07007_),
    .B1(_08793_),
    .Y(_08957_));
 sky130_fd_sc_hd__nor2_2 _36849_ (.A(_08956_),
    .B(_08957_),
    .Y(_08958_));
 sky130_fd_sc_hd__nor2_2 _36850_ (.A(_05504_),
    .B(_05440_),
    .Y(_08959_));
 sky130_fd_sc_hd__xor2_2 _36851_ (.A(_08958_),
    .B(_08959_),
    .X(_08960_));
 sky130_fd_sc_hd__nand2_2 _36852_ (.A(_00567_),
    .B(_07472_),
    .Y(_08961_));
 sky130_fd_sc_hd__nand2_2 _36853_ (.A(_00567_),
    .B(_07461_),
    .Y(_08963_));
 sky130_fd_sc_hd__o21ai_2 _36854_ (.A1(_07259_),
    .A2(_06023_),
    .B1(_08963_),
    .Y(_08964_));
 sky130_fd_sc_hd__o21ai_2 _36855_ (.A1(_08801_),
    .A2(_08961_),
    .B1(_08964_),
    .Y(_08965_));
 sky130_fd_sc_hd__nand2_2 _36856_ (.A(_06983_),
    .B(_08613_),
    .Y(_08966_));
 sky130_fd_sc_hd__xnor2_2 _36857_ (.A(_08965_),
    .B(_08966_),
    .Y(_08967_));
 sky130_fd_sc_hd__o22a_2 _36858_ (.A1(_08609_),
    .A2(_08963_),
    .B1(_08802_),
    .B2(_08803_),
    .X(_08968_));
 sky130_fd_sc_hd__xor2_2 _36859_ (.A(_08967_),
    .B(_08968_),
    .X(_08969_));
 sky130_fd_sc_hd__nand2_2 _36860_ (.A(_08960_),
    .B(_08969_),
    .Y(_08970_));
 sky130_fd_sc_hd__or2_2 _36861_ (.A(_08960_),
    .B(_08969_),
    .X(_08971_));
 sky130_fd_sc_hd__nand2_2 _36862_ (.A(_08970_),
    .B(_08971_),
    .Y(_08972_));
 sky130_fd_sc_hd__a21oi_2 _36863_ (.A1(_08806_),
    .A2(_08810_),
    .B1(_08972_),
    .Y(_08974_));
 sky130_fd_sc_hd__and3_2 _36864_ (.A(_08806_),
    .B(_08810_),
    .C(_08972_),
    .X(_08975_));
 sky130_fd_sc_hd__nor2_2 _36865_ (.A(_08974_),
    .B(_08975_),
    .Y(_08976_));
 sky130_fd_sc_hd__xnor2_2 _36866_ (.A(_08955_),
    .B(_08976_),
    .Y(_08977_));
 sky130_fd_sc_hd__or2_2 _36867_ (.A(_08954_),
    .B(_08977_),
    .X(_08978_));
 sky130_fd_sc_hd__nand2_2 _36868_ (.A(_08954_),
    .B(_08977_),
    .Y(_08979_));
 sky130_fd_sc_hd__and2_2 _36869_ (.A(_08978_),
    .B(_08979_),
    .X(_08980_));
 sky130_fd_sc_hd__o21a_2 _36870_ (.A1(_08788_),
    .A2(_08936_),
    .B1(_08980_),
    .X(_08981_));
 sky130_fd_sc_hd__nor3_2 _36871_ (.A(_08788_),
    .B(_08936_),
    .C(_08980_),
    .Y(_08982_));
 sky130_fd_sc_hd__nor2_2 _36872_ (.A(_08981_),
    .B(_08982_),
    .Y(_08983_));
 sky130_fd_sc_hd__xnor2_2 _36873_ (.A(_08935_),
    .B(_08983_),
    .Y(_08985_));
 sky130_fd_sc_hd__inv_2 _36874_ (.A(_08821_),
    .Y(_08986_));
 sky130_fd_sc_hd__nand2_2 _36875_ (.A(_08760_),
    .B(_08768_),
    .Y(_08987_));
 sky130_fd_sc_hd__o21ai_2 _36876_ (.A1(_08769_),
    .A2(_08986_),
    .B1(_08987_),
    .Y(_08988_));
 sky130_fd_sc_hd__xor2_2 _36877_ (.A(_08985_),
    .B(_08988_),
    .X(_08989_));
 sky130_fd_sc_hd__o21ba_2 _36878_ (.A1(_08791_),
    .A2(_08814_),
    .B1_N(_08813_),
    .X(_08990_));
 sky130_fd_sc_hd__xnor2_2 _36879_ (.A(_08818_),
    .B(_08990_),
    .Y(_08991_));
 sky130_fd_sc_hd__xnor2_2 _36880_ (.A(_08989_),
    .B(_08991_),
    .Y(_08992_));
 sky130_fd_sc_hd__or2b_2 _36881_ (.A(_08825_),
    .B_N(_08822_),
    .X(_08993_));
 sky130_fd_sc_hd__a21bo_2 _36882_ (.A1(_08826_),
    .A2(_08830_),
    .B1_N(_08993_),
    .X(_08994_));
 sky130_fd_sc_hd__xor2_2 _36883_ (.A(_08992_),
    .B(_08994_),
    .X(_08996_));
 sky130_fd_sc_hd__xor2_2 _36884_ (.A(_08828_),
    .B(_08996_),
    .X(_08997_));
 sky130_fd_sc_hd__o21a_2 _36885_ (.A1(_08922_),
    .A2(_08923_),
    .B1(_08997_),
    .X(_08998_));
 sky130_fd_sc_hd__inv_2 _36886_ (.A(_08998_),
    .Y(_08999_));
 sky130_fd_sc_hd__or3_2 _36887_ (.A(_08922_),
    .B(_08923_),
    .C(_08997_),
    .X(_09000_));
 sky130_fd_sc_hd__nand2_2 _36888_ (.A(_08999_),
    .B(_09000_),
    .Y(_09001_));
 sky130_fd_sc_hd__or2b_2 _36889_ (.A(_08648_),
    .B_N(_08838_),
    .X(_09002_));
 sky130_fd_sc_hd__a21oi_2 _36890_ (.A1(_08650_),
    .A2(_08655_),
    .B1(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__nor2_2 _36891_ (.A(_08836_),
    .B(_08837_),
    .Y(_09004_));
 sky130_fd_sc_hd__a21o_2 _36892_ (.A1(_08839_),
    .A2(_08838_),
    .B1(_09004_),
    .X(_09005_));
 sky130_fd_sc_hd__nor2_2 _36893_ (.A(_09003_),
    .B(_09005_),
    .Y(_09007_));
 sky130_fd_sc_hd__xnor2_2 _36894_ (.A(_09001_),
    .B(_09007_),
    .Y(_09008_));
 sky130_fd_sc_hd__and2b_2 _36895_ (.A_N(_08900_),
    .B(_08901_),
    .X(_09009_));
 sky130_fd_sc_hd__nand2_2 _36896_ (.A(iY[55]),
    .B(iX[63]),
    .Y(_09010_));
 sky130_fd_sc_hd__and2_2 _36897_ (.A(iY[57]),
    .B(iX[62]),
    .X(_09011_));
 sky130_fd_sc_hd__and3_2 _36898_ (.A(iY[56]),
    .B(iX[61]),
    .C(_09011_),
    .X(_09012_));
 sky130_fd_sc_hd__a22oi_2 _36899_ (.A1(iY[57]),
    .A2(iX[61]),
    .B1(iX[62]),
    .B2(iY[56]),
    .Y(_09013_));
 sky130_fd_sc_hd__o2bb2a_2 _36900_ (.A1_N(iY[58]),
    .A2_N(iX[60]),
    .B1(_09012_),
    .B2(_09013_),
    .X(_09014_));
 sky130_fd_sc_hd__and4bb_2 _36901_ (.A_N(_09012_),
    .B_N(_09013_),
    .C(iY[58]),
    .D(iX[60]),
    .X(_09015_));
 sky130_fd_sc_hd__nor2_2 _36902_ (.A(_09014_),
    .B(_09015_),
    .Y(_09016_));
 sky130_fd_sc_hd__xnor2_2 _36903_ (.A(_08845_),
    .B(_09016_),
    .Y(_09018_));
 sky130_fd_sc_hd__o21ai_2 _36904_ (.A1(_08850_),
    .A2(_08851_),
    .B1(_08848_),
    .Y(_09019_));
 sky130_fd_sc_hd__xor2_2 _36905_ (.A(_09018_),
    .B(_09019_),
    .X(_09020_));
 sky130_fd_sc_hd__a21bo_2 _36906_ (.A1(_08847_),
    .A2(_08852_),
    .B1_N(_08856_),
    .X(_09021_));
 sky130_fd_sc_hd__xor2_2 _36907_ (.A(_09020_),
    .B(_09021_),
    .X(_09022_));
 sky130_fd_sc_hd__xor2_2 _36908_ (.A(_08859_),
    .B(_09022_),
    .X(_09023_));
 sky130_fd_sc_hd__or2b_2 _36909_ (.A(_08874_),
    .B_N(_08873_),
    .X(_09024_));
 sky130_fd_sc_hd__and4_2 _36910_ (.A(iX[58]),
    .B(iX[59]),
    .C(iY[59]),
    .D(iY[60]),
    .X(_09025_));
 sky130_fd_sc_hd__a22oi_2 _36911_ (.A1(iX[59]),
    .A2(iY[59]),
    .B1(iY[60]),
    .B2(iX[58]),
    .Y(_09026_));
 sky130_fd_sc_hd__nor2_2 _36912_ (.A(_09025_),
    .B(_09026_),
    .Y(_09027_));
 sky130_fd_sc_hd__nand2_2 _36913_ (.A(iX[57]),
    .B(iY[61]),
    .Y(_09029_));
 sky130_fd_sc_hd__xnor2_2 _36914_ (.A(_09027_),
    .B(_09029_),
    .Y(_09030_));
 sky130_fd_sc_hd__o21ba_2 _36915_ (.A1(_08870_),
    .A2(_08872_),
    .B1_N(_08869_),
    .X(_09031_));
 sky130_fd_sc_hd__xnor2_2 _36916_ (.A(_09030_),
    .B(_09031_),
    .Y(_09032_));
 sky130_fd_sc_hd__and2_2 _36917_ (.A(iX[56]),
    .B(iY[62]),
    .X(_09033_));
 sky130_fd_sc_hd__or2_2 _36918_ (.A(_09032_),
    .B(_09033_),
    .X(_09034_));
 sky130_fd_sc_hd__nand2_2 _36919_ (.A(_09032_),
    .B(_09033_),
    .Y(_09035_));
 sky130_fd_sc_hd__nand2_2 _36920_ (.A(_09034_),
    .B(_09035_),
    .Y(_09036_));
 sky130_fd_sc_hd__a21oi_2 _36921_ (.A1(_09024_),
    .A2(_08879_),
    .B1(_09036_),
    .Y(_09037_));
 sky130_fd_sc_hd__and3_2 _36922_ (.A(_09024_),
    .B(_08879_),
    .C(_09036_),
    .X(_09038_));
 sky130_fd_sc_hd__nor2_2 _36923_ (.A(_09037_),
    .B(_09038_),
    .Y(_09040_));
 sky130_fd_sc_hd__nand2_2 _36924_ (.A(iX[55]),
    .B(iY[63]),
    .Y(_09041_));
 sky130_fd_sc_hd__xnor2_2 _36925_ (.A(_09040_),
    .B(_09041_),
    .Y(_09042_));
 sky130_fd_sc_hd__or2_2 _36926_ (.A(_09023_),
    .B(_09042_),
    .X(_09043_));
 sky130_fd_sc_hd__nand2_2 _36927_ (.A(_09023_),
    .B(_09042_),
    .Y(_09044_));
 sky130_fd_sc_hd__nand2_2 _36928_ (.A(_09043_),
    .B(_09044_),
    .Y(_09045_));
 sky130_fd_sc_hd__a21oi_2 _36929_ (.A1(_08867_),
    .A2(_08885_),
    .B1(_08865_),
    .Y(_09046_));
 sky130_fd_sc_hd__xnor2_2 _36930_ (.A(_09045_),
    .B(_09046_),
    .Y(_09047_));
 sky130_fd_sc_hd__nor2_2 _36931_ (.A(_09010_),
    .B(_09047_),
    .Y(_09048_));
 sky130_fd_sc_hd__and2_2 _36932_ (.A(_09010_),
    .B(_09047_),
    .X(_09049_));
 sky130_fd_sc_hd__nor2_2 _36933_ (.A(_09048_),
    .B(_09049_),
    .Y(_09051_));
 sky130_fd_sc_hd__o21ba_2 _36934_ (.A1(_08846_),
    .A2(_08890_),
    .B1_N(_08888_),
    .X(_09052_));
 sky130_fd_sc_hd__xnor2_2 _36935_ (.A(_09051_),
    .B(_09052_),
    .Y(_09053_));
 sky130_fd_sc_hd__o21ai_2 _36936_ (.A1(_08709_),
    .A2(_08895_),
    .B1(_08894_),
    .Y(_09054_));
 sky130_fd_sc_hd__nand2_2 _36937_ (.A(_09053_),
    .B(_09054_),
    .Y(_09055_));
 sky130_fd_sc_hd__or2_2 _36938_ (.A(_09053_),
    .B(_09054_),
    .X(_09056_));
 sky130_fd_sc_hd__nand2_2 _36939_ (.A(_09055_),
    .B(_09056_),
    .Y(_09057_));
 sky130_fd_sc_hd__a31o_2 _36940_ (.A1(iX[54]),
    .A2(iY[63]),
    .A3(_08883_),
    .B1(_08881_),
    .X(_09058_));
 sky130_fd_sc_hd__xnor2_2 _36941_ (.A(_09057_),
    .B(_09058_),
    .Y(_09059_));
 sky130_fd_sc_hd__o21ai_2 _36942_ (.A1(_08898_),
    .A2(_09009_),
    .B1(_09059_),
    .Y(_09060_));
 sky130_fd_sc_hd__or3_2 _36943_ (.A(_08898_),
    .B(_09009_),
    .C(_09059_),
    .X(_09062_));
 sky130_fd_sc_hd__and2_2 _36944_ (.A(_09060_),
    .B(_09062_),
    .X(_09063_));
 sky130_fd_sc_hd__a2111oi_2 _36945_ (.A1(_08732_),
    .A2(_08735_),
    .B1(_08904_),
    .C1(_08905_),
    .D1(_08730_),
    .Y(_09064_));
 sky130_fd_sc_hd__a21oi_2 _36946_ (.A1(_08728_),
    .A2(_08903_),
    .B1(_08905_),
    .Y(_09065_));
 sky130_fd_sc_hd__nor2_2 _36947_ (.A(_09064_),
    .B(_09065_),
    .Y(_09066_));
 sky130_fd_sc_hd__xnor2_2 _36948_ (.A(_09063_),
    .B(_09066_),
    .Y(_09067_));
 sky130_fd_sc_hd__xor2_2 _36949_ (.A(_09008_),
    .B(_09067_),
    .X(_09068_));
 sky130_fd_sc_hd__xnor2_2 _36950_ (.A(_17605_),
    .B(_09068_),
    .Y(_09069_));
 sky130_fd_sc_hd__inv_2 _36951_ (.A(_08909_),
    .Y(_09070_));
 sky130_fd_sc_hd__nand2_2 _36952_ (.A(_08841_),
    .B(_09070_),
    .Y(_09071_));
 sky130_fd_sc_hd__nand2_2 _36953_ (.A(_17259_),
    .B(_08910_),
    .Y(_09073_));
 sky130_fd_sc_hd__and2_2 _36954_ (.A(_09071_),
    .B(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__xnor2_2 _36955_ (.A(_09069_),
    .B(_09074_),
    .Y(_09075_));
 sky130_fd_sc_hd__a21oi_2 _36956_ (.A1(_08743_),
    .A2(_08913_),
    .B1(_08912_),
    .Y(_09076_));
 sky130_fd_sc_hd__inv_2 _36957_ (.A(_09076_),
    .Y(_09077_));
 sky130_fd_sc_hd__a31o_2 _36958_ (.A1(_08746_),
    .A2(_08749_),
    .A3(_08914_),
    .B1(_09077_),
    .X(_09078_));
 sky130_fd_sc_hd__xnor2_2 _36959_ (.A(_09075_),
    .B(_09078_),
    .Y(_09079_));
 sky130_fd_sc_hd__and2_2 _36960_ (.A(_17869_),
    .B(_09079_),
    .X(_09080_));
 sky130_fd_sc_hd__nor2_2 _36961_ (.A(_17869_),
    .B(_09079_),
    .Y(_09081_));
 sky130_fd_sc_hd__or2_2 _36962_ (.A(_09080_),
    .B(_09081_),
    .X(_09082_));
 sky130_fd_sc_hd__nand2_2 _36963_ (.A(_17376_),
    .B(_08916_),
    .Y(_09084_));
 sky130_fd_sc_hd__a21oi_2 _36964_ (.A1(_08751_),
    .A2(_09084_),
    .B1(_08918_),
    .Y(_09085_));
 sky130_fd_sc_hd__a21oi_2 _36965_ (.A1(_08754_),
    .A2(_08920_),
    .B1(_09085_),
    .Y(_09086_));
 sky130_fd_sc_hd__xor2_2 _36966_ (.A(_09082_),
    .B(_09086_),
    .X(oO[86]));
 sky130_fd_sc_hd__xor2_2 _36967_ (.A(_09069_),
    .B(_09074_),
    .X(_09087_));
 sky130_fd_sc_hd__a21o_2 _36968_ (.A1(_09071_),
    .A2(_09073_),
    .B1(_09069_),
    .X(_09088_));
 sky130_fd_sc_hd__a21bo_2 _36969_ (.A1(_09087_),
    .A2(_09078_),
    .B1_N(_09088_),
    .X(_09089_));
 sky130_fd_sc_hd__nor2_2 _36970_ (.A(_09008_),
    .B(_09067_),
    .Y(_09090_));
 sky130_fd_sc_hd__a21o_2 _36971_ (.A1(_17605_),
    .A2(_09068_),
    .B1(_09090_),
    .X(_09091_));
 sky130_fd_sc_hd__o21bai_2 _36972_ (.A1(_09003_),
    .A2(_09005_),
    .B1_N(_09001_),
    .Y(_09092_));
 sky130_fd_sc_hd__and2b_2 _36973_ (.A_N(_08992_),
    .B(_08994_),
    .X(_09094_));
 sky130_fd_sc_hd__nor2_2 _36974_ (.A(_08828_),
    .B(_08996_),
    .Y(_09095_));
 sky130_fd_sc_hd__and2b_2 _36975_ (.A_N(_08990_),
    .B(_08818_),
    .X(_09096_));
 sky130_fd_sc_hd__a21oi_2 _36976_ (.A1(_08958_),
    .A2(_08959_),
    .B1(_08956_),
    .Y(_09097_));
 sky130_fd_sc_hd__or2_2 _36977_ (.A(_08967_),
    .B(_08968_),
    .X(_09098_));
 sky130_fd_sc_hd__nor2_2 _36978_ (.A(_05227_),
    .B(_07252_),
    .Y(_09099_));
 sky130_fd_sc_hd__and3_2 _36979_ (.A(_06822_),
    .B(_04781_),
    .C(_09099_),
    .X(_09100_));
 sky130_fd_sc_hd__o22a_2 _36980_ (.A1(_05227_),
    .A2(_04782_),
    .B1(_08795_),
    .B2(_06816_),
    .X(_09101_));
 sky130_fd_sc_hd__nor2_2 _36981_ (.A(_09100_),
    .B(_09101_),
    .Y(_09102_));
 sky130_fd_sc_hd__nor2_2 _36982_ (.A(_05522_),
    .B(_05441_),
    .Y(_09103_));
 sky130_fd_sc_hd__xor2_2 _36983_ (.A(_09102_),
    .B(_09103_),
    .X(_09105_));
 sky130_fd_sc_hd__or3_2 _36984_ (.A(_07259_),
    .B(_08582_),
    .C(_08961_),
    .X(_09106_));
 sky130_fd_sc_hd__o21ai_2 _36985_ (.A1(_07259_),
    .A2(_08582_),
    .B1(_08961_),
    .Y(_09107_));
 sky130_fd_sc_hd__nand2_2 _36986_ (.A(_09106_),
    .B(_09107_),
    .Y(_09108_));
 sky130_fd_sc_hd__nand2_2 _36987_ (.A(_07461_),
    .B(_08613_),
    .Y(_09109_));
 sky130_fd_sc_hd__xnor2_2 _36988_ (.A(_09108_),
    .B(_09109_),
    .Y(_09110_));
 sky130_fd_sc_hd__o22a_2 _36989_ (.A1(_08801_),
    .A2(_08961_),
    .B1(_08965_),
    .B2(_08966_),
    .X(_09111_));
 sky130_fd_sc_hd__or2_2 _36990_ (.A(_09110_),
    .B(_09111_),
    .X(_09112_));
 sky130_fd_sc_hd__nand2_2 _36991_ (.A(_09110_),
    .B(_09111_),
    .Y(_09113_));
 sky130_fd_sc_hd__and2_2 _36992_ (.A(_09112_),
    .B(_09113_),
    .X(_09114_));
 sky130_fd_sc_hd__nand2_2 _36993_ (.A(_09105_),
    .B(_09114_),
    .Y(_09116_));
 sky130_fd_sc_hd__or2_2 _36994_ (.A(_09105_),
    .B(_09114_),
    .X(_09117_));
 sky130_fd_sc_hd__nand2_2 _36995_ (.A(_09116_),
    .B(_09117_),
    .Y(_09118_));
 sky130_fd_sc_hd__a21oi_2 _36996_ (.A1(_09098_),
    .A2(_08970_),
    .B1(_09118_),
    .Y(_09119_));
 sky130_fd_sc_hd__and3_2 _36997_ (.A(_09098_),
    .B(_08970_),
    .C(_09118_),
    .X(_09120_));
 sky130_fd_sc_hd__nor2_2 _36998_ (.A(_09119_),
    .B(_09120_),
    .Y(_09121_));
 sky130_fd_sc_hd__xnor2_2 _36999_ (.A(_09097_),
    .B(_09121_),
    .Y(_09122_));
 sky130_fd_sc_hd__inv_2 _37000_ (.A(_08948_),
    .Y(_09123_));
 sky130_fd_sc_hd__or2_2 _37001_ (.A(_08938_),
    .B(_08942_),
    .X(_09124_));
 sky130_fd_sc_hd__o22a_2 _37002_ (.A1(_03341_),
    .A2(_08571_),
    .B1(_08394_),
    .B2(_18344_),
    .X(_09125_));
 sky130_fd_sc_hd__a31oi_2 _37003_ (.A1(_07279_),
    .A2(_06783_),
    .A3(_08772_),
    .B1(_09125_),
    .Y(_09127_));
 sky130_fd_sc_hd__xnor2_2 _37004_ (.A(_09124_),
    .B(_09127_),
    .Y(_09128_));
 sky130_fd_sc_hd__nor2_2 _37005_ (.A(_09123_),
    .B(_09128_),
    .Y(_09129_));
 sky130_fd_sc_hd__and3_2 _37006_ (.A(_08945_),
    .B(_09123_),
    .C(_09128_),
    .X(_09130_));
 sky130_fd_sc_hd__nor2_2 _37007_ (.A(_08945_),
    .B(_09128_),
    .Y(_09131_));
 sky130_fd_sc_hd__nor3_2 _37008_ (.A(_09129_),
    .B(_09130_),
    .C(_09131_),
    .Y(_09132_));
 sky130_fd_sc_hd__and2_2 _37009_ (.A(_09122_),
    .B(_09132_),
    .X(_09133_));
 sky130_fd_sc_hd__nor2_2 _37010_ (.A(_09122_),
    .B(_09132_),
    .Y(_09134_));
 sky130_fd_sc_hd__or2_2 _37011_ (.A(_09133_),
    .B(_09134_),
    .X(_09135_));
 sky130_fd_sc_hd__a21oi_2 _37012_ (.A1(_08950_),
    .A2(_08978_),
    .B1(_09135_),
    .Y(_09136_));
 sky130_fd_sc_hd__and3_2 _37013_ (.A(_08950_),
    .B(_08978_),
    .C(_09135_),
    .X(_09138_));
 sky130_fd_sc_hd__nor2_2 _37014_ (.A(_09136_),
    .B(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__nor2_2 _37015_ (.A(_08926_),
    .B(_07533_),
    .Y(_09140_));
 sky130_fd_sc_hd__o22a_2 _37016_ (.A1(_05504_),
    .A2(_08931_),
    .B1(_08164_),
    .B2(_06491_),
    .X(_09141_));
 sky130_fd_sc_hd__nor2_2 _37017_ (.A(_09140_),
    .B(_09141_),
    .Y(_09142_));
 sky130_fd_sc_hd__o21ba_2 _37018_ (.A1(_08928_),
    .A2(_08932_),
    .B1_N(_08930_),
    .X(_09143_));
 sky130_fd_sc_hd__xnor2_2 _37019_ (.A(_09142_),
    .B(_09143_),
    .Y(_09144_));
 sky130_fd_sc_hd__xor2_2 _37020_ (.A(_09139_),
    .B(_09144_),
    .X(_09145_));
 sky130_fd_sc_hd__inv_2 _37021_ (.A(_08983_),
    .Y(_09146_));
 sky130_fd_sc_hd__nand2_2 _37022_ (.A(_08924_),
    .B(_08934_),
    .Y(_09147_));
 sky130_fd_sc_hd__o21ai_2 _37023_ (.A1(_08935_),
    .A2(_09146_),
    .B1(_09147_),
    .Y(_09149_));
 sky130_fd_sc_hd__xnor2_2 _37024_ (.A(_09145_),
    .B(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__a21oi_2 _37025_ (.A1(_08955_),
    .A2(_08976_),
    .B1(_08974_),
    .Y(_09151_));
 sky130_fd_sc_hd__xnor2_2 _37026_ (.A(_08981_),
    .B(_09151_),
    .Y(_09152_));
 sky130_fd_sc_hd__xnor2_2 _37027_ (.A(_09150_),
    .B(_09152_),
    .Y(_09153_));
 sky130_fd_sc_hd__nand2_2 _37028_ (.A(_08985_),
    .B(_08988_),
    .Y(_09154_));
 sky130_fd_sc_hd__a21boi_2 _37029_ (.A1(_08989_),
    .A2(_08991_),
    .B1_N(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__xnor2_2 _37030_ (.A(_09153_),
    .B(_09155_),
    .Y(_09156_));
 sky130_fd_sc_hd__xor2_2 _37031_ (.A(_09096_),
    .B(_09156_),
    .X(_09157_));
 sky130_fd_sc_hd__or3_2 _37032_ (.A(_09094_),
    .B(_09095_),
    .C(_09157_),
    .X(_09158_));
 sky130_fd_sc_hd__inv_2 _37033_ (.A(_09158_),
    .Y(_09160_));
 sky130_fd_sc_hd__o21a_2 _37034_ (.A1(_09094_),
    .A2(_09095_),
    .B1(_09157_),
    .X(_09161_));
 sky130_fd_sc_hd__nor2_2 _37035_ (.A(_09160_),
    .B(_09161_),
    .Y(_09162_));
 sky130_fd_sc_hd__a21o_2 _37036_ (.A1(_08999_),
    .A2(_09092_),
    .B1(_09162_),
    .X(_09163_));
 sky130_fd_sc_hd__nand3_2 _37037_ (.A(_08999_),
    .B(_09092_),
    .C(_09162_),
    .Y(_09164_));
 sky130_fd_sc_hd__or2b_2 _37038_ (.A(_09057_),
    .B_N(_09058_),
    .X(_09165_));
 sky130_fd_sc_hd__or2b_2 _37039_ (.A(_09052_),
    .B_N(_09051_),
    .X(_09166_));
 sky130_fd_sc_hd__and2b_2 _37040_ (.A_N(_09020_),
    .B(_09021_),
    .X(_09167_));
 sky130_fd_sc_hd__and3_2 _37041_ (.A(iY[56]),
    .B(iX[63]),
    .C(_09011_),
    .X(_09168_));
 sky130_fd_sc_hd__a21oi_2 _37042_ (.A1(iY[56]),
    .A2(iX[63]),
    .B1(_09011_),
    .Y(_09169_));
 sky130_fd_sc_hd__nand2_2 _37043_ (.A(iY[58]),
    .B(iX[61]),
    .Y(_09171_));
 sky130_fd_sc_hd__o21a_2 _37044_ (.A1(_09168_),
    .A2(_09169_),
    .B1(_09171_),
    .X(_09172_));
 sky130_fd_sc_hd__nor3_2 _37045_ (.A(_09168_),
    .B(_09169_),
    .C(_09171_),
    .Y(_09173_));
 sky130_fd_sc_hd__nor2_2 _37046_ (.A(_09172_),
    .B(_09173_),
    .Y(_09174_));
 sky130_fd_sc_hd__o21a_2 _37047_ (.A1(_09012_),
    .A2(_09015_),
    .B1(_09174_),
    .X(_09175_));
 sky130_fd_sc_hd__or3_2 _37048_ (.A(_09012_),
    .B(_09015_),
    .C(_09174_),
    .X(_09176_));
 sky130_fd_sc_hd__or2b_2 _37049_ (.A(_09175_),
    .B_N(_09176_),
    .X(_09177_));
 sky130_fd_sc_hd__and2b_2 _37050_ (.A_N(_09018_),
    .B(_09019_),
    .X(_09178_));
 sky130_fd_sc_hd__a21oi_2 _37051_ (.A1(_08845_),
    .A2(_09016_),
    .B1(_09178_),
    .Y(_09179_));
 sky130_fd_sc_hd__xor2_2 _37052_ (.A(_09177_),
    .B(_09179_),
    .X(_09180_));
 sky130_fd_sc_hd__xnor2_2 _37053_ (.A(_09167_),
    .B(_09180_),
    .Y(_09182_));
 sky130_fd_sc_hd__or2b_2 _37054_ (.A(_09031_),
    .B_N(_09030_),
    .X(_09183_));
 sky130_fd_sc_hd__and4_2 _37055_ (.A(iX[59]),
    .B(iY[59]),
    .C(iX[60]),
    .D(iY[60]),
    .X(_09184_));
 sky130_fd_sc_hd__a22oi_2 _37056_ (.A1(iY[59]),
    .A2(iX[60]),
    .B1(iY[60]),
    .B2(iX[59]),
    .Y(_09185_));
 sky130_fd_sc_hd__nor2_2 _37057_ (.A(_09184_),
    .B(_09185_),
    .Y(_09186_));
 sky130_fd_sc_hd__nand2_2 _37058_ (.A(iX[58]),
    .B(iY[61]),
    .Y(_09187_));
 sky130_fd_sc_hd__xnor2_2 _37059_ (.A(_09186_),
    .B(_09187_),
    .Y(_09188_));
 sky130_fd_sc_hd__o21ba_2 _37060_ (.A1(_09026_),
    .A2(_09029_),
    .B1_N(_09025_),
    .X(_09189_));
 sky130_fd_sc_hd__xnor2_2 _37061_ (.A(_09188_),
    .B(_09189_),
    .Y(_09190_));
 sky130_fd_sc_hd__and2_2 _37062_ (.A(iX[57]),
    .B(iY[62]),
    .X(_09191_));
 sky130_fd_sc_hd__or2_2 _37063_ (.A(_09190_),
    .B(_09191_),
    .X(_09193_));
 sky130_fd_sc_hd__nand2_2 _37064_ (.A(_09190_),
    .B(_09191_),
    .Y(_09194_));
 sky130_fd_sc_hd__nand2_2 _37065_ (.A(_09193_),
    .B(_09194_),
    .Y(_09195_));
 sky130_fd_sc_hd__a21oi_2 _37066_ (.A1(_09183_),
    .A2(_09035_),
    .B1(_09195_),
    .Y(_09196_));
 sky130_fd_sc_hd__and3_2 _37067_ (.A(_09183_),
    .B(_09035_),
    .C(_09195_),
    .X(_09197_));
 sky130_fd_sc_hd__nor2_2 _37068_ (.A(_09196_),
    .B(_09197_),
    .Y(_09198_));
 sky130_fd_sc_hd__nand2_2 _37069_ (.A(iX[56]),
    .B(iY[63]),
    .Y(_09199_));
 sky130_fd_sc_hd__xnor2_2 _37070_ (.A(_09198_),
    .B(_09199_),
    .Y(_09200_));
 sky130_fd_sc_hd__xnor2_2 _37071_ (.A(_09182_),
    .B(_09200_),
    .Y(_09201_));
 sky130_fd_sc_hd__o21ai_2 _37072_ (.A1(_08859_),
    .A2(_09022_),
    .B1(_09044_),
    .Y(_09202_));
 sky130_fd_sc_hd__and2_2 _37073_ (.A(_09201_),
    .B(_09202_),
    .X(_09204_));
 sky130_fd_sc_hd__nor2_2 _37074_ (.A(_09201_),
    .B(_09202_),
    .Y(_09205_));
 sky130_fd_sc_hd__nor2_2 _37075_ (.A(_09204_),
    .B(_09205_),
    .Y(_09206_));
 sky130_fd_sc_hd__o21bai_2 _37076_ (.A1(_09045_),
    .A2(_09046_),
    .B1_N(_09048_),
    .Y(_09207_));
 sky130_fd_sc_hd__xnor2_2 _37077_ (.A(_09206_),
    .B(_09207_),
    .Y(_09208_));
 sky130_fd_sc_hd__nor2_2 _37078_ (.A(_09166_),
    .B(_09208_),
    .Y(_09209_));
 sky130_fd_sc_hd__and2_2 _37079_ (.A(_09166_),
    .B(_09208_),
    .X(_09210_));
 sky130_fd_sc_hd__nor2_2 _37080_ (.A(_09209_),
    .B(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__a31o_2 _37081_ (.A1(iX[55]),
    .A2(iY[63]),
    .A3(_09040_),
    .B1(_09037_),
    .X(_09212_));
 sky130_fd_sc_hd__xnor2_2 _37082_ (.A(_09211_),
    .B(_09212_),
    .Y(_09213_));
 sky130_fd_sc_hd__a21oi_2 _37083_ (.A1(_09055_),
    .A2(_09165_),
    .B1(_09213_),
    .Y(_09215_));
 sky130_fd_sc_hd__and3_2 _37084_ (.A(_09055_),
    .B(_09165_),
    .C(_09213_),
    .X(_09216_));
 sky130_fd_sc_hd__nor2_2 _37085_ (.A(_09215_),
    .B(_09216_),
    .Y(_09217_));
 sky130_fd_sc_hd__inv_2 _37086_ (.A(_09063_),
    .Y(_09218_));
 sky130_fd_sc_hd__o21a_2 _37087_ (.A1(_09218_),
    .A2(_09066_),
    .B1(_09060_),
    .X(_09219_));
 sky130_fd_sc_hd__xnor2_2 _37088_ (.A(_09217_),
    .B(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__nand3_2 _37089_ (.A(_09163_),
    .B(_09164_),
    .C(_09220_),
    .Y(_09221_));
 sky130_fd_sc_hd__a21o_2 _37090_ (.A1(_09163_),
    .A2(_09164_),
    .B1(_09220_),
    .X(_09222_));
 sky130_fd_sc_hd__nand3_2 _37091_ (.A(_17944_),
    .B(_09221_),
    .C(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__a21o_2 _37092_ (.A1(_09221_),
    .A2(_09222_),
    .B1(_17944_),
    .X(_09224_));
 sky130_fd_sc_hd__and2_2 _37093_ (.A(_09223_),
    .B(_09224_),
    .X(_09226_));
 sky130_fd_sc_hd__buf_1 _37094_ (.A(_09226_),
    .X(_09227_));
 sky130_fd_sc_hd__xor2_2 _37095_ (.A(_09091_),
    .B(_09227_),
    .X(_09228_));
 sky130_fd_sc_hd__xnor2_2 _37096_ (.A(_09089_),
    .B(_09228_),
    .Y(_09229_));
 sky130_fd_sc_hd__nor2_2 _37097_ (.A(_18080_),
    .B(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__nand2_2 _37098_ (.A(_18080_),
    .B(_09229_),
    .Y(_09231_));
 sky130_fd_sc_hd__and2b_2 _37099_ (.A_N(_09230_),
    .B(_09231_),
    .X(_09232_));
 sky130_fd_sc_hd__o21ba_2 _37100_ (.A1(_09082_),
    .A2(_09086_),
    .B1_N(_09080_),
    .X(_09233_));
 sky130_fd_sc_hd__xnor2_2 _37101_ (.A(_09232_),
    .B(_09233_),
    .Y(oO[87]));
 sky130_fd_sc_hd__nor3b_2 _37102_ (.A(_09082_),
    .B(_09230_),
    .C_N(_09231_),
    .Y(_09234_));
 sky130_fd_sc_hd__and3_2 _37103_ (.A(_08753_),
    .B(_08920_),
    .C(_09234_),
    .X(_09236_));
 sky130_fd_sc_hd__nand4_2 _37104_ (.A(_07932_),
    .B(_08158_),
    .C(_08556_),
    .D(_09236_),
    .Y(_09237_));
 sky130_fd_sc_hd__a21bo_2 _37105_ (.A1(_08363_),
    .A2(_08556_),
    .B1_N(_08558_),
    .X(_09238_));
 sky130_fd_sc_hd__a221o_2 _37106_ (.A1(_09080_),
    .A2(_09231_),
    .B1(_09234_),
    .B2(_09085_),
    .C1(_09230_),
    .X(_09239_));
 sky130_fd_sc_hd__a21o_2 _37107_ (.A1(_09236_),
    .A2(_09238_),
    .B1(_09239_),
    .X(_09240_));
 sky130_fd_sc_hd__o21ba_2 _37108_ (.A1(_07945_),
    .A2(_09237_),
    .B1_N(_09240_),
    .X(_09241_));
 sky130_fd_sc_hd__and2b_2 _37109_ (.A_N(_09151_),
    .B(_08981_),
    .X(_09242_));
 sky130_fd_sc_hd__nand2_2 _37110_ (.A(_09145_),
    .B(_09149_),
    .Y(_09243_));
 sky130_fd_sc_hd__inv_2 _37111_ (.A(_09243_),
    .Y(_09244_));
 sky130_fd_sc_hd__or2_2 _37112_ (.A(_09145_),
    .B(_09149_),
    .X(_09245_));
 sky130_fd_sc_hd__and3_2 _37113_ (.A(_09243_),
    .B(_09245_),
    .C(_09152_),
    .X(_09247_));
 sky130_fd_sc_hd__nand2_2 _37114_ (.A(_09139_),
    .B(_09144_),
    .Y(_09248_));
 sky130_fd_sc_hd__a21oi_2 _37115_ (.A1(_08930_),
    .A2(_09142_),
    .B1(_09140_),
    .Y(_09249_));
 sky130_fd_sc_hd__nand2_2 _37116_ (.A(_08933_),
    .B(_09142_),
    .Y(_09250_));
 sky130_fd_sc_hd__a311o_2 _37117_ (.A1(_08561_),
    .A2(_08925_),
    .A3(_08927_),
    .B1(_09250_),
    .C1(_08764_),
    .X(_09251_));
 sky130_fd_sc_hd__nor2_2 _37118_ (.A(_08926_),
    .B(_07534_),
    .Y(_09252_));
 sky130_fd_sc_hd__o22a_2 _37119_ (.A1(_05522_),
    .A2(_08931_),
    .B1(_08164_),
    .B2(_18344_),
    .X(_09253_));
 sky130_fd_sc_hd__or2_2 _37120_ (.A(_09252_),
    .B(_09253_),
    .X(_09254_));
 sky130_fd_sc_hd__a21o_2 _37121_ (.A1(_09249_),
    .A2(_09251_),
    .B1(_09254_),
    .X(_09255_));
 sky130_fd_sc_hd__nand3_2 _37122_ (.A(_09254_),
    .B(_09249_),
    .C(_09251_),
    .Y(_09256_));
 sky130_fd_sc_hd__a21oi_2 _37123_ (.A1(_09102_),
    .A2(_09103_),
    .B1(_09100_),
    .Y(_09258_));
 sky130_fd_sc_hd__nand2_2 _37124_ (.A(_07461_),
    .B(_07007_),
    .Y(_09259_));
 sky130_fd_sc_hd__xnor2_2 _37125_ (.A(_09099_),
    .B(_09259_),
    .Y(_09260_));
 sky130_fd_sc_hd__nor2_2 _37126_ (.A(_06816_),
    .B(_07983_),
    .Y(_09261_));
 sky130_fd_sc_hd__xor2_2 _37127_ (.A(_09260_),
    .B(_09261_),
    .X(_09262_));
 sky130_fd_sc_hd__nor2_2 _37128_ (.A(_07259_),
    .B(_08582_),
    .Y(_09263_));
 sky130_fd_sc_hd__nor2_2 _37129_ (.A(_02311_),
    .B(_06797_),
    .Y(_09264_));
 sky130_fd_sc_hd__o22a_2 _37130_ (.A1(_02311_),
    .A2(_08582_),
    .B1(_08571_),
    .B2(_07259_),
    .X(_09265_));
 sky130_fd_sc_hd__a21o_2 _37131_ (.A1(_09263_),
    .A2(_09264_),
    .B1(_09265_),
    .X(_09266_));
 sky130_fd_sc_hd__nand2_2 _37132_ (.A(_08613_),
    .B(_07472_),
    .Y(_09267_));
 sky130_fd_sc_hd__xnor2_2 _37133_ (.A(_09266_),
    .B(_09267_),
    .Y(_09269_));
 sky130_fd_sc_hd__o21a_2 _37134_ (.A1(_09108_),
    .A2(_09109_),
    .B1(_09106_),
    .X(_09270_));
 sky130_fd_sc_hd__or2_2 _37135_ (.A(_09269_),
    .B(_09270_),
    .X(_09271_));
 sky130_fd_sc_hd__nand2_2 _37136_ (.A(_09269_),
    .B(_09270_),
    .Y(_09272_));
 sky130_fd_sc_hd__and2_2 _37137_ (.A(_09271_),
    .B(_09272_),
    .X(_09273_));
 sky130_fd_sc_hd__nand2_2 _37138_ (.A(_09262_),
    .B(_09273_),
    .Y(_09274_));
 sky130_fd_sc_hd__or2_2 _37139_ (.A(_09262_),
    .B(_09273_),
    .X(_09275_));
 sky130_fd_sc_hd__nand2_2 _37140_ (.A(_09274_),
    .B(_09275_),
    .Y(_09276_));
 sky130_fd_sc_hd__a21oi_2 _37141_ (.A1(_09112_),
    .A2(_09116_),
    .B1(_09276_),
    .Y(_09277_));
 sky130_fd_sc_hd__and3_2 _37142_ (.A(_09112_),
    .B(_09116_),
    .C(_09276_),
    .X(_09278_));
 sky130_fd_sc_hd__nor2_2 _37143_ (.A(_09277_),
    .B(_09278_),
    .Y(_09280_));
 sky130_fd_sc_hd__xnor2_2 _37144_ (.A(_09258_),
    .B(_09280_),
    .Y(_09281_));
 sky130_fd_sc_hd__o211a_2 _37145_ (.A1(_18344_),
    .A2(_08571_),
    .B1(_06783_),
    .C1(_07279_),
    .X(_09282_));
 sky130_fd_sc_hd__and2_2 _37146_ (.A(_09124_),
    .B(_09127_),
    .X(_09283_));
 sky130_fd_sc_hd__nor2_2 _37147_ (.A(_09283_),
    .B(_09131_),
    .Y(_09284_));
 sky130_fd_sc_hd__xnor2_2 _37148_ (.A(_09282_),
    .B(_09284_),
    .Y(_09285_));
 sky130_fd_sc_hd__and2_2 _37149_ (.A(_09281_),
    .B(_09285_),
    .X(_09286_));
 sky130_fd_sc_hd__nor2_2 _37150_ (.A(_09281_),
    .B(_09285_),
    .Y(_09287_));
 sky130_fd_sc_hd__nor2_2 _37151_ (.A(_09286_),
    .B(_09287_),
    .Y(_09288_));
 sky130_fd_sc_hd__o21a_2 _37152_ (.A1(_09129_),
    .A2(_09133_),
    .B1(_09288_),
    .X(_09289_));
 sky130_fd_sc_hd__nor3_2 _37153_ (.A(_09129_),
    .B(_09133_),
    .C(_09288_),
    .Y(_09291_));
 sky130_fd_sc_hd__nor2_2 _37154_ (.A(_09289_),
    .B(_09291_),
    .Y(_09292_));
 sky130_fd_sc_hd__and3_2 _37155_ (.A(_09255_),
    .B(_09256_),
    .C(_09292_),
    .X(_09293_));
 sky130_fd_sc_hd__a21oi_2 _37156_ (.A1(_09255_),
    .A2(_09256_),
    .B1(_09292_),
    .Y(_09294_));
 sky130_fd_sc_hd__or3_2 _37157_ (.A(_09248_),
    .B(_09293_),
    .C(_09294_),
    .X(_09295_));
 sky130_fd_sc_hd__o21ai_2 _37158_ (.A1(_09293_),
    .A2(_09294_),
    .B1(_09248_),
    .Y(_09296_));
 sky130_fd_sc_hd__o21ba_2 _37159_ (.A1(_09097_),
    .A2(_09120_),
    .B1_N(_09119_),
    .X(_09297_));
 sky130_fd_sc_hd__xnor2_2 _37160_ (.A(_09136_),
    .B(_09297_),
    .Y(_09298_));
 sky130_fd_sc_hd__nand3_2 _37161_ (.A(_09295_),
    .B(_09296_),
    .C(_09298_),
    .Y(_09299_));
 sky130_fd_sc_hd__a21o_2 _37162_ (.A1(_09295_),
    .A2(_09296_),
    .B1(_09298_),
    .X(_09300_));
 sky130_fd_sc_hd__o211ai_2 _37163_ (.A1(_09244_),
    .A2(_09247_),
    .B1(_09299_),
    .C1(_09300_),
    .Y(_09302_));
 sky130_fd_sc_hd__a211o_2 _37164_ (.A1(_09299_),
    .A2(_09300_),
    .B1(_09244_),
    .C1(_09247_),
    .X(_09303_));
 sky130_fd_sc_hd__and3_2 _37165_ (.A(_09242_),
    .B(_09302_),
    .C(_09303_),
    .X(_09304_));
 sky130_fd_sc_hd__a21oi_2 _37166_ (.A1(_09302_),
    .A2(_09303_),
    .B1(_09242_),
    .Y(_09305_));
 sky130_fd_sc_hd__nor2_2 _37167_ (.A(_09304_),
    .B(_09305_),
    .Y(_09306_));
 sky130_fd_sc_hd__and2_2 _37168_ (.A(_09243_),
    .B(_09245_),
    .X(_09307_));
 sky130_fd_sc_hd__nor2_2 _37169_ (.A(_09307_),
    .B(_09152_),
    .Y(_09308_));
 sky130_fd_sc_hd__nand2_2 _37170_ (.A(_09096_),
    .B(_09156_),
    .Y(_09309_));
 sky130_fd_sc_hd__o31ai_2 _37171_ (.A1(_09247_),
    .A2(_09308_),
    .A3(_09155_),
    .B1(_09309_),
    .Y(_09310_));
 sky130_fd_sc_hd__xnor2_2 _37172_ (.A(_09306_),
    .B(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__a21o_2 _37173_ (.A1(_08650_),
    .A2(_08655_),
    .B1(_09002_),
    .X(_09313_));
 sky130_fd_sc_hd__o21a_2 _37174_ (.A1(_08998_),
    .A2(_09161_),
    .B1(_09158_),
    .X(_09314_));
 sky130_fd_sc_hd__nor2_2 _37175_ (.A(_09005_),
    .B(_09314_),
    .Y(_09315_));
 sky130_fd_sc_hd__o21a_2 _37176_ (.A1(_09000_),
    .A2(_09161_),
    .B1(_09158_),
    .X(_09316_));
 sky130_fd_sc_hd__inv_2 _37177_ (.A(_09316_),
    .Y(_09317_));
 sky130_fd_sc_hd__a21oi_2 _37178_ (.A1(_09313_),
    .A2(_09315_),
    .B1(_09317_),
    .Y(_09318_));
 sky130_fd_sc_hd__xnor2_2 _37179_ (.A(_09311_),
    .B(_09318_),
    .Y(_09319_));
 sky130_fd_sc_hd__nor2_2 _37180_ (.A(_09060_),
    .B(_09216_),
    .Y(_09320_));
 sky130_fd_sc_hd__or3_2 _37181_ (.A(_09065_),
    .B(_09215_),
    .C(_09320_),
    .X(_09321_));
 sky130_fd_sc_hd__inv_2 _37182_ (.A(_09216_),
    .Y(_09322_));
 sky130_fd_sc_hd__a21o_2 _37183_ (.A1(_09062_),
    .A2(_09322_),
    .B1(_09215_),
    .X(_09324_));
 sky130_fd_sc_hd__a31o_2 _37184_ (.A1(iX[56]),
    .A2(iY[63]),
    .A3(_09198_),
    .B1(_09196_),
    .X(_09325_));
 sky130_fd_sc_hd__or2b_2 _37185_ (.A(_09189_),
    .B_N(_09188_),
    .X(_09326_));
 sky130_fd_sc_hd__and4_2 _37186_ (.A(iY[59]),
    .B(iX[60]),
    .C(iY[60]),
    .D(iX[61]),
    .X(_09327_));
 sky130_fd_sc_hd__a22oi_2 _37187_ (.A1(iX[60]),
    .A2(iY[60]),
    .B1(iX[61]),
    .B2(iY[59]),
    .Y(_09328_));
 sky130_fd_sc_hd__nor2_2 _37188_ (.A(_09327_),
    .B(_09328_),
    .Y(_09329_));
 sky130_fd_sc_hd__nand2_2 _37189_ (.A(iX[59]),
    .B(iY[61]),
    .Y(_09330_));
 sky130_fd_sc_hd__xnor2_2 _37190_ (.A(_09329_),
    .B(_09330_),
    .Y(_09331_));
 sky130_fd_sc_hd__o21ba_2 _37191_ (.A1(_09185_),
    .A2(_09187_),
    .B1_N(_09184_),
    .X(_09332_));
 sky130_fd_sc_hd__xnor2_2 _37192_ (.A(_09331_),
    .B(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__and2_2 _37193_ (.A(iX[58]),
    .B(iY[62]),
    .X(_09335_));
 sky130_fd_sc_hd__or2_2 _37194_ (.A(_09333_),
    .B(_09335_),
    .X(_09336_));
 sky130_fd_sc_hd__nand2_2 _37195_ (.A(_09333_),
    .B(_09335_),
    .Y(_09337_));
 sky130_fd_sc_hd__nand2_2 _37196_ (.A(_09336_),
    .B(_09337_),
    .Y(_09338_));
 sky130_fd_sc_hd__a21oi_2 _37197_ (.A1(_09326_),
    .A2(_09194_),
    .B1(_09338_),
    .Y(_09339_));
 sky130_fd_sc_hd__and3_2 _37198_ (.A(_09326_),
    .B(_09194_),
    .C(_09338_),
    .X(_09340_));
 sky130_fd_sc_hd__nor2_2 _37199_ (.A(_09339_),
    .B(_09340_),
    .Y(_09341_));
 sky130_fd_sc_hd__nand2_2 _37200_ (.A(iX[57]),
    .B(iY[63]),
    .Y(_09342_));
 sky130_fd_sc_hd__xnor2_2 _37201_ (.A(_09341_),
    .B(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__nor2_2 _37202_ (.A(_09177_),
    .B(_09179_),
    .Y(_09344_));
 sky130_fd_sc_hd__nand2_2 _37203_ (.A(iY[57]),
    .B(iX[62]),
    .Y(_09346_));
 sky130_fd_sc_hd__nand2_2 _37204_ (.A(iY[58]),
    .B(iX[63]),
    .Y(_09347_));
 sky130_fd_sc_hd__a22o_2 _37205_ (.A1(iY[58]),
    .A2(iX[62]),
    .B1(iX[63]),
    .B2(iY[57]),
    .X(_09348_));
 sky130_fd_sc_hd__o21a_2 _37206_ (.A1(_09346_),
    .A2(_09347_),
    .B1(_09348_),
    .X(_09349_));
 sky130_fd_sc_hd__o21ai_2 _37207_ (.A1(_09168_),
    .A2(_09173_),
    .B1(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__or3_2 _37208_ (.A(_09168_),
    .B(_09173_),
    .C(_09349_),
    .X(_09351_));
 sky130_fd_sc_hd__and2_2 _37209_ (.A(_09350_),
    .B(_09351_),
    .X(_09352_));
 sky130_fd_sc_hd__nand2_2 _37210_ (.A(_09344_),
    .B(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__or3_2 _37211_ (.A(_09175_),
    .B(_09344_),
    .C(_09352_),
    .X(_09354_));
 sky130_fd_sc_hd__nand2_2 _37212_ (.A(_09175_),
    .B(_09352_),
    .Y(_09355_));
 sky130_fd_sc_hd__and3_2 _37213_ (.A(_09353_),
    .B(_09354_),
    .C(_09355_),
    .X(_09357_));
 sky130_fd_sc_hd__xnor2_2 _37214_ (.A(_09343_),
    .B(_09357_),
    .Y(_09358_));
 sky130_fd_sc_hd__and2b_2 _37215_ (.A_N(_09182_),
    .B(_09200_),
    .X(_09359_));
 sky130_fd_sc_hd__a21o_2 _37216_ (.A1(_09167_),
    .A2(_09180_),
    .B1(_09359_),
    .X(_09360_));
 sky130_fd_sc_hd__and2b_2 _37217_ (.A_N(_09358_),
    .B(_09360_),
    .X(_09361_));
 sky130_fd_sc_hd__and2b_2 _37218_ (.A_N(_09360_),
    .B(_09358_),
    .X(_09362_));
 sky130_fd_sc_hd__nor2_2 _37219_ (.A(_09361_),
    .B(_09362_),
    .Y(_09363_));
 sky130_fd_sc_hd__a21o_2 _37220_ (.A1(_09206_),
    .A2(_09207_),
    .B1(_09204_),
    .X(_09364_));
 sky130_fd_sc_hd__xnor2_2 _37221_ (.A(_09363_),
    .B(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__xor2_2 _37222_ (.A(_09325_),
    .B(_09365_),
    .X(_09366_));
 sky130_fd_sc_hd__a21oi_2 _37223_ (.A1(_09211_),
    .A2(_09212_),
    .B1(_09209_),
    .Y(_09368_));
 sky130_fd_sc_hd__nor2_2 _37224_ (.A(_09366_),
    .B(_09368_),
    .Y(_09369_));
 sky130_fd_sc_hd__and2_2 _37225_ (.A(_09366_),
    .B(_09368_),
    .X(_09370_));
 sky130_fd_sc_hd__nor2_2 _37226_ (.A(_09369_),
    .B(_09370_),
    .Y(_09371_));
 sky130_fd_sc_hd__o211a_2 _37227_ (.A1(_09064_),
    .A2(_09321_),
    .B1(_09324_),
    .C1(_09371_),
    .X(_09372_));
 sky130_fd_sc_hd__o21a_2 _37228_ (.A1(_09064_),
    .A2(_09321_),
    .B1(_09324_),
    .X(_09373_));
 sky130_fd_sc_hd__nor2_2 _37229_ (.A(_09371_),
    .B(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__nor2_2 _37230_ (.A(_09372_),
    .B(_09374_),
    .Y(_09375_));
 sky130_fd_sc_hd__xnor2_2 _37231_ (.A(_09319_),
    .B(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__and2_2 _37232_ (.A(_18312_),
    .B(_09376_),
    .X(_09377_));
 sky130_fd_sc_hd__nor2_2 _37233_ (.A(_18312_),
    .B(_09376_),
    .Y(_09379_));
 sky130_fd_sc_hd__or2_2 _37234_ (.A(_09377_),
    .B(_09379_),
    .X(_09380_));
 sky130_fd_sc_hd__and2_2 _37235_ (.A(_09222_),
    .B(_09223_),
    .X(_09381_));
 sky130_fd_sc_hd__or2_2 _37236_ (.A(_09380_),
    .B(_09381_),
    .X(_09382_));
 sky130_fd_sc_hd__nand2_2 _37237_ (.A(_09380_),
    .B(_09381_),
    .Y(_09383_));
 sky130_fd_sc_hd__and2_2 _37238_ (.A(_09382_),
    .B(_09383_),
    .X(_09384_));
 sky130_fd_sc_hd__and3_2 _37239_ (.A(_08746_),
    .B(_09087_),
    .C(_09228_),
    .X(_09385_));
 sky130_fd_sc_hd__nor2_2 _37240_ (.A(_09091_),
    .B(_09227_),
    .Y(_09386_));
 sky130_fd_sc_hd__nand2_2 _37241_ (.A(_09091_),
    .B(_09227_),
    .Y(_09387_));
 sky130_fd_sc_hd__o21bai_2 _37242_ (.A1(_09091_),
    .A2(_09227_),
    .B1_N(_09088_),
    .Y(_09388_));
 sky130_fd_sc_hd__o311ai_2 _37243_ (.A1(_09075_),
    .A2(_09076_),
    .A3(_09386_),
    .B1(_09387_),
    .C1(_09388_),
    .Y(_09390_));
 sky130_fd_sc_hd__a31o_4 _37244_ (.A1(_08749_),
    .A2(_08914_),
    .A3(_09385_),
    .B1(_09390_),
    .X(_09391_));
 sky130_fd_sc_hd__xor2_2 _37245_ (.A(_09384_),
    .B(_09391_),
    .X(_09392_));
 sky130_fd_sc_hd__and2_2 _37246_ (.A(_18647_),
    .B(_09392_),
    .X(_09393_));
 sky130_fd_sc_hd__nor2_2 _37247_ (.A(_18647_),
    .B(_09392_),
    .Y(_09394_));
 sky130_fd_sc_hd__nor2_2 _37248_ (.A(_09393_),
    .B(_09394_),
    .Y(_09395_));
 sky130_fd_sc_hd__and2b_2 _37249_ (.A_N(_09241_),
    .B(_09395_),
    .X(_09396_));
 sky130_fd_sc_hd__and2b_2 _37250_ (.A_N(_09395_),
    .B(_09241_),
    .X(_09397_));
 sky130_fd_sc_hd__nor2_2 _37251_ (.A(_09396_),
    .B(_09397_),
    .Y(oO[88]));
 sky130_fd_sc_hd__and2b_2 _37252_ (.A_N(_09297_),
    .B(_09136_),
    .X(_09398_));
 sky130_fd_sc_hd__and2_2 _37253_ (.A(_09131_),
    .B(_09282_),
    .X(_09400_));
 sky130_fd_sc_hd__and3_2 _37254_ (.A(_07461_),
    .B(_07007_),
    .C(_09099_),
    .X(_09401_));
 sky130_fd_sc_hd__a21o_2 _37255_ (.A1(_09260_),
    .A2(_09261_),
    .B1(_09401_),
    .X(_09402_));
 sky130_fd_sc_hd__or3_2 _37256_ (.A(_06023_),
    .B(_08795_),
    .C(_09259_),
    .X(_09403_));
 sky130_fd_sc_hd__a2bb2o_2 _37257_ (.A1_N(_05543_),
    .A2_N(_08795_),
    .B1(_07007_),
    .B2(_07472_),
    .X(_09404_));
 sky130_fd_sc_hd__nand2_2 _37258_ (.A(_09403_),
    .B(_09404_),
    .Y(_09405_));
 sky130_fd_sc_hd__nor2_2 _37259_ (.A(_05227_),
    .B(_07983_),
    .Y(_09406_));
 sky130_fd_sc_hd__xnor2_2 _37260_ (.A(_09405_),
    .B(_09406_),
    .Y(_09407_));
 sky130_fd_sc_hd__nor2_2 _37261_ (.A(_07259_),
    .B(_05550_),
    .Y(_09408_));
 sky130_fd_sc_hd__xnor2_2 _37262_ (.A(_09264_),
    .B(_09408_),
    .Y(_09409_));
 sky130_fd_sc_hd__nand2_2 _37263_ (.A(_08613_),
    .B(_06154_),
    .Y(_09411_));
 sky130_fd_sc_hd__nor2_2 _37264_ (.A(_09409_),
    .B(_09411_),
    .Y(_09412_));
 sky130_fd_sc_hd__and2_2 _37265_ (.A(_09409_),
    .B(_09411_),
    .X(_09413_));
 sky130_fd_sc_hd__or2_2 _37266_ (.A(_09412_),
    .B(_09413_),
    .X(_09414_));
 sky130_fd_sc_hd__o2bb2a_2 _37267_ (.A1_N(_09263_),
    .A2_N(_09264_),
    .B1(_09265_),
    .B2(_09267_),
    .X(_09415_));
 sky130_fd_sc_hd__or2_2 _37268_ (.A(_09414_),
    .B(_09415_),
    .X(_09416_));
 sky130_fd_sc_hd__nand2_2 _37269_ (.A(_09414_),
    .B(_09415_),
    .Y(_09417_));
 sky130_fd_sc_hd__and2_2 _37270_ (.A(_09416_),
    .B(_09417_),
    .X(_09418_));
 sky130_fd_sc_hd__nand2_2 _37271_ (.A(_09407_),
    .B(_09418_),
    .Y(_09419_));
 sky130_fd_sc_hd__or2_2 _37272_ (.A(_09407_),
    .B(_09418_),
    .X(_09420_));
 sky130_fd_sc_hd__nand2_2 _37273_ (.A(_09419_),
    .B(_09420_),
    .Y(_09422_));
 sky130_fd_sc_hd__a21oi_2 _37274_ (.A1(_09271_),
    .A2(_09274_),
    .B1(_09422_),
    .Y(_09423_));
 sky130_fd_sc_hd__and3_2 _37275_ (.A(_09271_),
    .B(_09274_),
    .C(_09422_),
    .X(_09424_));
 sky130_fd_sc_hd__nor2_2 _37276_ (.A(_09423_),
    .B(_09424_),
    .Y(_09425_));
 sky130_fd_sc_hd__xor2_2 _37277_ (.A(_09402_),
    .B(_09425_),
    .X(_09426_));
 sky130_fd_sc_hd__o211a_2 _37278_ (.A1(_08772_),
    .A2(_09283_),
    .B1(_07279_),
    .C1(_06783_),
    .X(_09427_));
 sky130_fd_sc_hd__and2_2 _37279_ (.A(_09426_),
    .B(_09427_),
    .X(_09428_));
 sky130_fd_sc_hd__nor2_2 _37280_ (.A(_09426_),
    .B(_09427_),
    .Y(_09429_));
 sky130_fd_sc_hd__nor2_2 _37281_ (.A(_09428_),
    .B(_09429_),
    .Y(_09430_));
 sky130_fd_sc_hd__o21a_2 _37282_ (.A1(_09286_),
    .A2(_09400_),
    .B1(_09430_),
    .X(_09431_));
 sky130_fd_sc_hd__nor3_2 _37283_ (.A(_09286_),
    .B(_09430_),
    .C(_09400_),
    .Y(_09433_));
 sky130_fd_sc_hd__nor2_2 _37284_ (.A(_09431_),
    .B(_09433_),
    .Y(_09434_));
 sky130_fd_sc_hd__o22a_2 _37285_ (.A1(_06816_),
    .A2(_08931_),
    .B1(_08164_),
    .B2(_03341_),
    .X(_09435_));
 sky130_fd_sc_hd__and3_2 _37286_ (.A(_07279_),
    .B(_06822_),
    .C(_08763_),
    .X(_09436_));
 sky130_fd_sc_hd__nor2_2 _37287_ (.A(_09435_),
    .B(_09436_),
    .Y(_09437_));
 sky130_fd_sc_hd__a21oi_2 _37288_ (.A1(_09249_),
    .A2(_09251_),
    .B1(_09254_),
    .Y(_09438_));
 sky130_fd_sc_hd__nor2_2 _37289_ (.A(_09252_),
    .B(_09438_),
    .Y(_09439_));
 sky130_fd_sc_hd__xnor2_2 _37290_ (.A(_09437_),
    .B(_09439_),
    .Y(_09440_));
 sky130_fd_sc_hd__xor2_2 _37291_ (.A(_09434_),
    .B(_09440_),
    .X(_09441_));
 sky130_fd_sc_hd__xnor2_2 _37292_ (.A(_09293_),
    .B(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__and2b_2 _37293_ (.A_N(_09258_),
    .B(_09280_),
    .X(_09444_));
 sky130_fd_sc_hd__o21a_2 _37294_ (.A1(_09277_),
    .A2(_09444_),
    .B1(_09289_),
    .X(_09445_));
 sky130_fd_sc_hd__nor3_2 _37295_ (.A(_09277_),
    .B(_09444_),
    .C(_09289_),
    .Y(_09446_));
 sky130_fd_sc_hd__or2_2 _37296_ (.A(_09445_),
    .B(_09446_),
    .X(_09447_));
 sky130_fd_sc_hd__nor2_2 _37297_ (.A(_09442_),
    .B(_09447_),
    .Y(_09448_));
 sky130_fd_sc_hd__and2_2 _37298_ (.A(_09442_),
    .B(_09447_),
    .X(_09449_));
 sky130_fd_sc_hd__a211o_2 _37299_ (.A1(_09295_),
    .A2(_09299_),
    .B1(_09448_),
    .C1(_09449_),
    .X(_09450_));
 sky130_fd_sc_hd__o211ai_2 _37300_ (.A1(_09448_),
    .A2(_09449_),
    .B1(_09295_),
    .C1(_09299_),
    .Y(_09451_));
 sky130_fd_sc_hd__and3_2 _37301_ (.A(_09398_),
    .B(_09450_),
    .C(_09451_),
    .X(_09452_));
 sky130_fd_sc_hd__a21oi_2 _37302_ (.A1(_09450_),
    .A2(_09451_),
    .B1(_09398_),
    .Y(_09453_));
 sky130_fd_sc_hd__nor2_2 _37303_ (.A(_09452_),
    .B(_09453_),
    .Y(_09455_));
 sky130_fd_sc_hd__a21bo_2 _37304_ (.A1(_09242_),
    .A2(_09303_),
    .B1_N(_09302_),
    .X(_09456_));
 sky130_fd_sc_hd__xnor2_2 _37305_ (.A(_09455_),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__or2_2 _37306_ (.A(_09306_),
    .B(_09310_),
    .X(_09458_));
 sky130_fd_sc_hd__nand2_2 _37307_ (.A(_09306_),
    .B(_09310_),
    .Y(_09459_));
 sky130_fd_sc_hd__a21bo_2 _37308_ (.A1(_09458_),
    .A2(_09318_),
    .B1_N(_09459_),
    .X(_09460_));
 sky130_fd_sc_hd__xnor2_2 _37309_ (.A(_09457_),
    .B(_09460_),
    .Y(_09461_));
 sky130_fd_sc_hd__and2b_2 _37310_ (.A_N(_09365_),
    .B(_09325_),
    .X(_09462_));
 sky130_fd_sc_hd__a31o_2 _37311_ (.A1(iX[57]),
    .A2(iY[63]),
    .A3(_09341_),
    .B1(_09339_),
    .X(_09463_));
 sky130_fd_sc_hd__or2b_2 _37312_ (.A(_09332_),
    .B_N(_09331_),
    .X(_09464_));
 sky130_fd_sc_hd__and4_2 _37313_ (.A(iY[59]),
    .B(iY[60]),
    .C(iX[61]),
    .D(iX[62]),
    .X(_09466_));
 sky130_fd_sc_hd__a22oi_2 _37314_ (.A1(iY[60]),
    .A2(iX[61]),
    .B1(iX[62]),
    .B2(iY[59]),
    .Y(_09467_));
 sky130_fd_sc_hd__nor2_2 _37315_ (.A(_09466_),
    .B(_09467_),
    .Y(_09468_));
 sky130_fd_sc_hd__nand2_2 _37316_ (.A(iX[60]),
    .B(iY[61]),
    .Y(_09469_));
 sky130_fd_sc_hd__xnor2_2 _37317_ (.A(_09468_),
    .B(_09469_),
    .Y(_09470_));
 sky130_fd_sc_hd__o21ba_2 _37318_ (.A1(_09328_),
    .A2(_09330_),
    .B1_N(_09327_),
    .X(_09471_));
 sky130_fd_sc_hd__xnor2_2 _37319_ (.A(_09470_),
    .B(_09471_),
    .Y(_09472_));
 sky130_fd_sc_hd__and2_2 _37320_ (.A(iX[59]),
    .B(iY[62]),
    .X(_09473_));
 sky130_fd_sc_hd__or2_2 _37321_ (.A(_09472_),
    .B(_09473_),
    .X(_09474_));
 sky130_fd_sc_hd__nand2_2 _37322_ (.A(_09472_),
    .B(_09473_),
    .Y(_09475_));
 sky130_fd_sc_hd__nand2_2 _37323_ (.A(_09474_),
    .B(_09475_),
    .Y(_09477_));
 sky130_fd_sc_hd__a21oi_2 _37324_ (.A1(_09464_),
    .A2(_09337_),
    .B1(_09477_),
    .Y(_09478_));
 sky130_fd_sc_hd__and3_2 _37325_ (.A(_09464_),
    .B(_09337_),
    .C(_09477_),
    .X(_09479_));
 sky130_fd_sc_hd__nor2_2 _37326_ (.A(_09478_),
    .B(_09479_),
    .Y(_09480_));
 sky130_fd_sc_hd__nand2_2 _37327_ (.A(iX[58]),
    .B(iY[63]),
    .Y(_09481_));
 sky130_fd_sc_hd__xnor2_2 _37328_ (.A(_09480_),
    .B(_09481_),
    .Y(_09482_));
 sky130_fd_sc_hd__and4b_2 _37329_ (.A_N(_09347_),
    .B(_09350_),
    .C(_09355_),
    .D(_09346_),
    .X(_09483_));
 sky130_fd_sc_hd__o2bb2a_2 _37330_ (.A1_N(_09350_),
    .A2_N(_09355_),
    .B1(_09011_),
    .B2(_09347_),
    .X(_09484_));
 sky130_fd_sc_hd__or2_2 _37331_ (.A(_09483_),
    .B(_09484_),
    .X(_09485_));
 sky130_fd_sc_hd__nand2_2 _37332_ (.A(_09482_),
    .B(_09485_),
    .Y(_09486_));
 sky130_fd_sc_hd__or2_2 _37333_ (.A(_09482_),
    .B(_09485_),
    .X(_09488_));
 sky130_fd_sc_hd__and2_2 _37334_ (.A(_09486_),
    .B(_09488_),
    .X(_09489_));
 sky130_fd_sc_hd__a22o_2 _37335_ (.A1(_09344_),
    .A2(_09352_),
    .B1(_09357_),
    .B2(_09343_),
    .X(_09490_));
 sky130_fd_sc_hd__and2_2 _37336_ (.A(_09489_),
    .B(_09490_),
    .X(_09491_));
 sky130_fd_sc_hd__nor2_2 _37337_ (.A(_09489_),
    .B(_09490_),
    .Y(_09492_));
 sky130_fd_sc_hd__nor2_2 _37338_ (.A(_09491_),
    .B(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__nand2_2 _37339_ (.A(_09361_),
    .B(_09493_),
    .Y(_09494_));
 sky130_fd_sc_hd__and3_2 _37340_ (.A(_09201_),
    .B(_09202_),
    .C(_09363_),
    .X(_09495_));
 sky130_fd_sc_hd__nand2_2 _37341_ (.A(_09493_),
    .B(_09495_),
    .Y(_09496_));
 sky130_fd_sc_hd__or3_2 _37342_ (.A(_09361_),
    .B(_09493_),
    .C(_09495_),
    .X(_09497_));
 sky130_fd_sc_hd__and3_2 _37343_ (.A(_09494_),
    .B(_09496_),
    .C(_09497_),
    .X(_09499_));
 sky130_fd_sc_hd__xor2_2 _37344_ (.A(_09463_),
    .B(_09499_),
    .X(_09500_));
 sky130_fd_sc_hd__and3_2 _37345_ (.A(_09206_),
    .B(_09207_),
    .C(_09363_),
    .X(_09501_));
 sky130_fd_sc_hd__nor3_2 _37346_ (.A(_09462_),
    .B(_09500_),
    .C(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__inv_2 _37347_ (.A(_09502_),
    .Y(_09503_));
 sky130_fd_sc_hd__o21ai_2 _37348_ (.A1(_09462_),
    .A2(_09501_),
    .B1(_09500_),
    .Y(_09504_));
 sky130_fd_sc_hd__nand2_2 _37349_ (.A(_09503_),
    .B(_09504_),
    .Y(_09505_));
 sky130_fd_sc_hd__nor2_2 _37350_ (.A(_09369_),
    .B(_09372_),
    .Y(_09506_));
 sky130_fd_sc_hd__xnor2_2 _37351_ (.A(_09505_),
    .B(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__xor2_2 _37352_ (.A(_09461_),
    .B(_09507_),
    .X(_09508_));
 sky130_fd_sc_hd__nand2_2 _37353_ (.A(_18714_),
    .B(_09508_),
    .Y(_09510_));
 sky130_fd_sc_hd__or2_2 _37354_ (.A(_18714_),
    .B(_09508_),
    .X(_09511_));
 sky130_fd_sc_hd__nand2_2 _37355_ (.A(_09510_),
    .B(_09511_),
    .Y(_09512_));
 sky130_fd_sc_hd__inv_2 _37356_ (.A(_09375_),
    .Y(_09513_));
 sky130_fd_sc_hd__a21oi_2 _37357_ (.A1(_09319_),
    .A2(_09513_),
    .B1(_09377_),
    .Y(_09514_));
 sky130_fd_sc_hd__nor2_2 _37358_ (.A(_09512_),
    .B(_09514_),
    .Y(_09515_));
 sky130_fd_sc_hd__and2_2 _37359_ (.A(_09512_),
    .B(_09514_),
    .X(_09516_));
 sky130_fd_sc_hd__nor2_2 _37360_ (.A(_09515_),
    .B(_09516_),
    .Y(_09517_));
 sky130_fd_sc_hd__a21boi_2 _37361_ (.A1(_09384_),
    .A2(_09391_),
    .B1_N(_09382_),
    .Y(_09518_));
 sky130_fd_sc_hd__xnor2_2 _37362_ (.A(_09517_),
    .B(_09518_),
    .Y(_09519_));
 sky130_fd_sc_hd__nor2_2 _37363_ (.A(_00076_),
    .B(_09519_),
    .Y(_09521_));
 sky130_fd_sc_hd__and2_2 _37364_ (.A(_00076_),
    .B(_09519_),
    .X(_09522_));
 sky130_fd_sc_hd__nor2_2 _37365_ (.A(_09521_),
    .B(_09522_),
    .Y(_09523_));
 sky130_fd_sc_hd__nor2_2 _37366_ (.A(_09393_),
    .B(_09396_),
    .Y(_09524_));
 sky130_fd_sc_hd__xnor2_2 _37367_ (.A(_09523_),
    .B(_09524_),
    .Y(oO[89]));
 sky130_fd_sc_hd__nand2_2 _37368_ (.A(_09461_),
    .B(_09507_),
    .Y(_09525_));
 sky130_fd_sc_hd__nand2_2 _37369_ (.A(_09434_),
    .B(_09440_),
    .Y(_09526_));
 sky130_fd_sc_hd__o22a_2 _37370_ (.A1(_05227_),
    .A2(_08931_),
    .B1(_08164_),
    .B2(_07259_),
    .X(_09527_));
 sky130_fd_sc_hd__a31o_2 _37371_ (.A1(_05450_),
    .A2(_06983_),
    .A3(_08763_),
    .B1(_09527_),
    .X(_09528_));
 sky130_fd_sc_hd__inv_2 _37372_ (.A(_09528_),
    .Y(_09529_));
 sky130_fd_sc_hd__inv_2 _37373_ (.A(_09435_),
    .Y(_09531_));
 sky130_fd_sc_hd__o311a_2 _37374_ (.A1(_09252_),
    .A2(_09438_),
    .A3(_09436_),
    .B1(_09529_),
    .C1(_09531_),
    .X(_09532_));
 sky130_fd_sc_hd__o31a_2 _37375_ (.A1(_09252_),
    .A2(_09438_),
    .A3(_09436_),
    .B1(_09531_),
    .X(_09533_));
 sky130_fd_sc_hd__nor2_2 _37376_ (.A(_09529_),
    .B(_09533_),
    .Y(_09534_));
 sky130_fd_sc_hd__or2_2 _37377_ (.A(_09532_),
    .B(_09534_),
    .X(_09535_));
 sky130_fd_sc_hd__o22a_2 _37378_ (.A1(_00944_),
    .A2(_08571_),
    .B1(_08394_),
    .B2(_02311_),
    .X(_09536_));
 sky130_fd_sc_hd__a31o_2 _37379_ (.A1(_08613_),
    .A2(_06783_),
    .A3(_09264_),
    .B1(_09536_),
    .X(_09537_));
 sky130_fd_sc_hd__a21oi_2 _37380_ (.A1(_09264_),
    .A2(_09408_),
    .B1(_09412_),
    .Y(_09538_));
 sky130_fd_sc_hd__nor2_2 _37381_ (.A(_09537_),
    .B(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__and2_2 _37382_ (.A(_09537_),
    .B(_09538_),
    .X(_09540_));
 sky130_fd_sc_hd__nor2_2 _37383_ (.A(_09539_),
    .B(_09540_),
    .Y(_09541_));
 sky130_fd_sc_hd__or4_2 _37384_ (.A(_06023_),
    .B(_04782_),
    .C(_08582_),
    .D(_08795_),
    .X(_09542_));
 sky130_fd_sc_hd__a2bb2o_2 _37385_ (.A1_N(_06023_),
    .A2_N(_08795_),
    .B1(_06154_),
    .B2(_07007_),
    .X(_09543_));
 sky130_fd_sc_hd__nand2_2 _37386_ (.A(_09542_),
    .B(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__nor2_2 _37387_ (.A(_05543_),
    .B(_07983_),
    .Y(_09545_));
 sky130_fd_sc_hd__xnor2_2 _37388_ (.A(_09544_),
    .B(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__xnor2_2 _37389_ (.A(_09541_),
    .B(_09546_),
    .Y(_09547_));
 sky130_fd_sc_hd__a21oi_2 _37390_ (.A1(_09416_),
    .A2(_09419_),
    .B1(_09547_),
    .Y(_09548_));
 sky130_fd_sc_hd__and3_2 _37391_ (.A(_09416_),
    .B(_09419_),
    .C(_09547_),
    .X(_09549_));
 sky130_fd_sc_hd__nor2_2 _37392_ (.A(_09548_),
    .B(_09549_),
    .Y(_09550_));
 sky130_fd_sc_hd__a21bo_2 _37393_ (.A1(_09404_),
    .A2(_09406_),
    .B1_N(_09403_),
    .X(_09552_));
 sky130_fd_sc_hd__xor2_2 _37394_ (.A(_09550_),
    .B(_09552_),
    .X(_09553_));
 sky130_fd_sc_hd__nand2_2 _37395_ (.A(_09428_),
    .B(_09553_),
    .Y(_09554_));
 sky130_fd_sc_hd__or2_2 _37396_ (.A(_09428_),
    .B(_09553_),
    .X(_09555_));
 sky130_fd_sc_hd__nand2_2 _37397_ (.A(_09554_),
    .B(_09555_),
    .Y(_09556_));
 sky130_fd_sc_hd__xor2_2 _37398_ (.A(_09535_),
    .B(_09556_),
    .X(_09557_));
 sky130_fd_sc_hd__xor2_2 _37399_ (.A(_09526_),
    .B(_09557_),
    .X(_09558_));
 sky130_fd_sc_hd__and2_2 _37400_ (.A(_09402_),
    .B(_09425_),
    .X(_09559_));
 sky130_fd_sc_hd__o21ai_2 _37401_ (.A1(_09423_),
    .A2(_09559_),
    .B1(_09431_),
    .Y(_09560_));
 sky130_fd_sc_hd__or3_2 _37402_ (.A(_09423_),
    .B(_09559_),
    .C(_09431_),
    .X(_09561_));
 sky130_fd_sc_hd__nand2_2 _37403_ (.A(_09560_),
    .B(_09561_),
    .Y(_09563_));
 sky130_fd_sc_hd__xor2_2 _37404_ (.A(_09558_),
    .B(_09563_),
    .X(_09564_));
 sky130_fd_sc_hd__a21oi_2 _37405_ (.A1(_09293_),
    .A2(_09441_),
    .B1(_09448_),
    .Y(_09565_));
 sky130_fd_sc_hd__xnor2_2 _37406_ (.A(_09564_),
    .B(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__xnor2_2 _37407_ (.A(_09445_),
    .B(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__inv_2 _37408_ (.A(_09450_),
    .Y(_09568_));
 sky130_fd_sc_hd__nor2_2 _37409_ (.A(_09568_),
    .B(_09452_),
    .Y(_09569_));
 sky130_fd_sc_hd__nor2_2 _37410_ (.A(_09567_),
    .B(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__nand2_2 _37411_ (.A(_09567_),
    .B(_09569_),
    .Y(_09571_));
 sky130_fd_sc_hd__or2b_2 _37412_ (.A(_09570_),
    .B_N(_09571_),
    .X(_09572_));
 sky130_fd_sc_hd__a2111o_2 _37413_ (.A1(_09313_),
    .A2(_09315_),
    .B1(_09317_),
    .C1(_09457_),
    .D1(_09311_),
    .X(_09574_));
 sky130_fd_sc_hd__nand2_2 _37414_ (.A(_09455_),
    .B(_09456_),
    .Y(_09575_));
 sky130_fd_sc_hd__o21a_2 _37415_ (.A1(_09459_),
    .A2(_09457_),
    .B1(_09575_),
    .X(_09576_));
 sky130_fd_sc_hd__and2_2 _37416_ (.A(_09574_),
    .B(_09576_),
    .X(_09577_));
 sky130_fd_sc_hd__xnor2_2 _37417_ (.A(_09572_),
    .B(_09577_),
    .Y(_09578_));
 sky130_fd_sc_hd__or3_2 _37418_ (.A(_09011_),
    .B(_09347_),
    .C(_09355_),
    .X(_09579_));
 sky130_fd_sc_hd__a21oi_2 _37419_ (.A1(_09346_),
    .A2(_09350_),
    .B1(_09347_),
    .Y(_09580_));
 sky130_fd_sc_hd__or2b_2 _37420_ (.A(_09471_),
    .B_N(_09470_),
    .X(_09581_));
 sky130_fd_sc_hd__nand2_2 _37421_ (.A(iY[60]),
    .B(iX[62]),
    .Y(_09582_));
 sky130_fd_sc_hd__nand2_2 _37422_ (.A(iY[59]),
    .B(iX[63]),
    .Y(_09583_));
 sky130_fd_sc_hd__and4_2 _37423_ (.A(iY[59]),
    .B(iY[60]),
    .C(iX[62]),
    .D(iX[63]),
    .X(_09585_));
 sky130_fd_sc_hd__a21o_2 _37424_ (.A1(_09582_),
    .A2(_09583_),
    .B1(_09585_),
    .X(_09586_));
 sky130_fd_sc_hd__nand2_2 _37425_ (.A(iX[61]),
    .B(iY[61]),
    .Y(_09587_));
 sky130_fd_sc_hd__xor2_2 _37426_ (.A(_09586_),
    .B(_09587_),
    .X(_09588_));
 sky130_fd_sc_hd__o21ba_2 _37427_ (.A1(_09467_),
    .A2(_09469_),
    .B1_N(_09466_),
    .X(_09589_));
 sky130_fd_sc_hd__xnor2_2 _37428_ (.A(_09588_),
    .B(_09589_),
    .Y(_09590_));
 sky130_fd_sc_hd__nand2_2 _37429_ (.A(iX[60]),
    .B(iY[62]),
    .Y(_09591_));
 sky130_fd_sc_hd__xor2_2 _37430_ (.A(_09590_),
    .B(_09591_),
    .X(_09592_));
 sky130_fd_sc_hd__a21oi_2 _37431_ (.A1(_09581_),
    .A2(_09475_),
    .B1(_09592_),
    .Y(_09593_));
 sky130_fd_sc_hd__and3_2 _37432_ (.A(_09581_),
    .B(_09475_),
    .C(_09592_),
    .X(_09594_));
 sky130_fd_sc_hd__nor2_2 _37433_ (.A(_09593_),
    .B(_09594_),
    .Y(_09596_));
 sky130_fd_sc_hd__nand2_2 _37434_ (.A(iX[59]),
    .B(iY[63]),
    .Y(_09597_));
 sky130_fd_sc_hd__xnor2_2 _37435_ (.A(_09596_),
    .B(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__xnor2_2 _37436_ (.A(_09580_),
    .B(_09598_),
    .Y(_09599_));
 sky130_fd_sc_hd__a21oi_2 _37437_ (.A1(_09579_),
    .A2(_09486_),
    .B1(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__and3_2 _37438_ (.A(_09579_),
    .B(_09486_),
    .C(_09599_),
    .X(_09601_));
 sky130_fd_sc_hd__nor2_2 _37439_ (.A(_09600_),
    .B(_09601_),
    .Y(_09602_));
 sky130_fd_sc_hd__nand2_2 _37440_ (.A(_09491_),
    .B(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__or2_2 _37441_ (.A(_09491_),
    .B(_09602_),
    .X(_09604_));
 sky130_fd_sc_hd__nand2_2 _37442_ (.A(_09603_),
    .B(_09604_),
    .Y(_09605_));
 sky130_fd_sc_hd__nor2_2 _37443_ (.A(_09494_),
    .B(_09605_),
    .Y(_09607_));
 sky130_fd_sc_hd__and2_2 _37444_ (.A(_09494_),
    .B(_09605_),
    .X(_09608_));
 sky130_fd_sc_hd__or2_2 _37445_ (.A(_09607_),
    .B(_09608_),
    .X(_09609_));
 sky130_fd_sc_hd__a31o_2 _37446_ (.A1(iX[58]),
    .A2(iY[63]),
    .A3(_09480_),
    .B1(_09478_),
    .X(_09610_));
 sky130_fd_sc_hd__xnor2_2 _37447_ (.A(_09609_),
    .B(_09610_),
    .Y(_09611_));
 sky130_fd_sc_hd__a22o_2 _37448_ (.A1(_09493_),
    .A2(_09495_),
    .B1(_09499_),
    .B2(_09463_),
    .X(_09612_));
 sky130_fd_sc_hd__and2_2 _37449_ (.A(_09611_),
    .B(_09612_),
    .X(_09613_));
 sky130_fd_sc_hd__nor2_2 _37450_ (.A(_09611_),
    .B(_09612_),
    .Y(_09614_));
 sky130_fd_sc_hd__nor2_2 _37451_ (.A(_09613_),
    .B(_09614_),
    .Y(_09615_));
 sky130_fd_sc_hd__inv_2 _37452_ (.A(_09504_),
    .Y(_09616_));
 sky130_fd_sc_hd__o31a_2 _37453_ (.A1(_09369_),
    .A2(_09372_),
    .A3(_09616_),
    .B1(_09503_),
    .X(_09618_));
 sky130_fd_sc_hd__and2_2 _37454_ (.A(_09615_),
    .B(_09618_),
    .X(_09619_));
 sky130_fd_sc_hd__nor2_2 _37455_ (.A(_09615_),
    .B(_09618_),
    .Y(_09620_));
 sky130_fd_sc_hd__nor2_2 _37456_ (.A(_09619_),
    .B(_09620_),
    .Y(_09621_));
 sky130_fd_sc_hd__xor2_2 _37457_ (.A(_09578_),
    .B(_09621_),
    .X(_09622_));
 sky130_fd_sc_hd__nand2b_2 _37458_ (.A_N(_00138_),
    .B(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__or2b_2 _37459_ (.A(_09622_),
    .B_N(_00138_),
    .X(_09624_));
 sky130_fd_sc_hd__nand2_2 _37460_ (.A(_09623_),
    .B(_09624_),
    .Y(_09625_));
 sky130_fd_sc_hd__a21oi_2 _37461_ (.A1(_09525_),
    .A2(_09510_),
    .B1(_09625_),
    .Y(_09626_));
 sky130_fd_sc_hd__and3_2 _37462_ (.A(_09525_),
    .B(_09510_),
    .C(_09625_),
    .X(_09627_));
 sky130_fd_sc_hd__nor2_2 _37463_ (.A(_09626_),
    .B(_09627_),
    .Y(_09629_));
 sky130_fd_sc_hd__or2_2 _37464_ (.A(_09512_),
    .B(_09514_),
    .X(_09630_));
 sky130_fd_sc_hd__a21oi_2 _37465_ (.A1(_09382_),
    .A2(_09630_),
    .B1(_09516_),
    .Y(_09631_));
 sky130_fd_sc_hd__a31o_2 _37466_ (.A1(_09384_),
    .A2(_09391_),
    .A3(_09517_),
    .B1(_09631_),
    .X(_09632_));
 sky130_fd_sc_hd__xor2_2 _37467_ (.A(_09629_),
    .B(_09632_),
    .X(_09633_));
 sky130_fd_sc_hd__and2_2 _37468_ (.A(_00469_),
    .B(_09633_),
    .X(_09634_));
 sky130_fd_sc_hd__nor2_2 _37469_ (.A(_00469_),
    .B(_09633_),
    .Y(_09635_));
 sky130_fd_sc_hd__nor2_2 _37470_ (.A(_09634_),
    .B(_09635_),
    .Y(_09636_));
 sky130_fd_sc_hd__or2_2 _37471_ (.A(_00076_),
    .B(_09519_),
    .X(_09637_));
 sky130_fd_sc_hd__o21a_2 _37472_ (.A1(_09393_),
    .A2(_09522_),
    .B1(_09637_),
    .X(_09638_));
 sky130_fd_sc_hd__a21o_2 _37473_ (.A1(_09396_),
    .A2(_09523_),
    .B1(_09638_),
    .X(_09640_));
 sky130_fd_sc_hd__xor2_2 _37474_ (.A(_09636_),
    .B(_09640_),
    .X(oO[90]));
 sky130_fd_sc_hd__a21o_2 _37475_ (.A1(_09629_),
    .A2(_09632_),
    .B1(_09626_),
    .X(_09641_));
 sky130_fd_sc_hd__or2_2 _37476_ (.A(_09578_),
    .B(_09621_),
    .X(_09642_));
 sky130_fd_sc_hd__and2b_2 _37477_ (.A_N(_09609_),
    .B(_09610_),
    .X(_09643_));
 sky130_fd_sc_hd__nor2_2 _37478_ (.A(_09586_),
    .B(_09587_),
    .Y(_09644_));
 sky130_fd_sc_hd__nand2_2 _37479_ (.A(iY[61]),
    .B(iX[63]),
    .Y(_09645_));
 sky130_fd_sc_hd__a22o_2 _37480_ (.A1(iY[61]),
    .A2(iX[62]),
    .B1(iX[63]),
    .B2(iY[60]),
    .X(_09646_));
 sky130_fd_sc_hd__o21a_2 _37481_ (.A1(_09582_),
    .A2(_09645_),
    .B1(_09646_),
    .X(_09647_));
 sky130_fd_sc_hd__o21a_2 _37482_ (.A1(_09585_),
    .A2(_09644_),
    .B1(_09647_),
    .X(_09648_));
 sky130_fd_sc_hd__nor3_2 _37483_ (.A(_09585_),
    .B(_09644_),
    .C(_09647_),
    .Y(_09650_));
 sky130_fd_sc_hd__nor2_2 _37484_ (.A(_09648_),
    .B(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__nand2_2 _37485_ (.A(iX[61]),
    .B(iY[62]),
    .Y(_09652_));
 sky130_fd_sc_hd__xor2_2 _37486_ (.A(_09651_),
    .B(_09652_),
    .X(_09653_));
 sky130_fd_sc_hd__and2b_2 _37487_ (.A_N(_09589_),
    .B(_09588_),
    .X(_09654_));
 sky130_fd_sc_hd__a31oi_2 _37488_ (.A1(iX[60]),
    .A2(iY[62]),
    .A3(_09590_),
    .B1(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__xnor2_2 _37489_ (.A(_09653_),
    .B(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__nand2_2 _37490_ (.A(iX[60]),
    .B(iY[63]),
    .Y(_09657_));
 sky130_fd_sc_hd__nor2_2 _37491_ (.A(_09656_),
    .B(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__and2_2 _37492_ (.A(_09656_),
    .B(_09657_),
    .X(_09659_));
 sky130_fd_sc_hd__nor2_2 _37493_ (.A(_09658_),
    .B(_09659_),
    .Y(_09661_));
 sky130_fd_sc_hd__a21oi_2 _37494_ (.A1(_09580_),
    .A2(_09598_),
    .B1(_09600_),
    .Y(_09662_));
 sky130_fd_sc_hd__xnor2_2 _37495_ (.A(_09661_),
    .B(_09662_),
    .Y(_09663_));
 sky130_fd_sc_hd__xnor2_2 _37496_ (.A(_09603_),
    .B(_09663_),
    .Y(_09664_));
 sky130_fd_sc_hd__o21ba_2 _37497_ (.A1(_09594_),
    .A2(_09597_),
    .B1_N(_09593_),
    .X(_09665_));
 sky130_fd_sc_hd__xnor2_2 _37498_ (.A(_09664_),
    .B(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__o21a_2 _37499_ (.A1(_09607_),
    .A2(_09643_),
    .B1(_09666_),
    .X(_09667_));
 sky130_fd_sc_hd__or3_2 _37500_ (.A(_09607_),
    .B(_09643_),
    .C(_09666_),
    .X(_09668_));
 sky130_fd_sc_hd__or2b_2 _37501_ (.A(_09667_),
    .B_N(_09668_),
    .X(_09669_));
 sky130_fd_sc_hd__or2_2 _37502_ (.A(_09613_),
    .B(_09619_),
    .X(_09670_));
 sky130_fd_sc_hd__xnor2_2 _37503_ (.A(_09669_),
    .B(_09670_),
    .Y(_09672_));
 sky130_fd_sc_hd__and3_2 _37504_ (.A(_09434_),
    .B(_09440_),
    .C(_09557_),
    .X(_09673_));
 sky130_fd_sc_hd__nor2_2 _37505_ (.A(_09558_),
    .B(_09563_),
    .Y(_09674_));
 sky130_fd_sc_hd__nor2_2 _37506_ (.A(_09535_),
    .B(_09556_),
    .Y(_09675_));
 sky130_fd_sc_hd__a21bo_2 _37507_ (.A1(_09543_),
    .A2(_09545_),
    .B1_N(_09542_),
    .X(_09676_));
 sky130_fd_sc_hd__nor2_2 _37508_ (.A(_08795_),
    .B(_08571_),
    .Y(_09677_));
 sky130_fd_sc_hd__and3_2 _37509_ (.A(_07007_),
    .B(_06154_),
    .C(_09677_),
    .X(_09678_));
 sky130_fd_sc_hd__o22a_2 _37510_ (.A1(_08582_),
    .A2(_08795_),
    .B1(_08571_),
    .B2(_04782_),
    .X(_09679_));
 sky130_fd_sc_hd__nor2_2 _37511_ (.A(_09678_),
    .B(_09679_),
    .Y(_09680_));
 sky130_fd_sc_hd__nor2_2 _37512_ (.A(_06023_),
    .B(_07983_),
    .Y(_09681_));
 sky130_fd_sc_hd__xor2_2 _37513_ (.A(_09680_),
    .B(_09681_),
    .X(_09683_));
 sky130_fd_sc_hd__or3_2 _37514_ (.A(_00944_),
    .B(_08394_),
    .C(_09264_),
    .X(_09684_));
 sky130_fd_sc_hd__xor2_2 _37515_ (.A(_09683_),
    .B(_09684_),
    .X(_09685_));
 sky130_fd_sc_hd__a21o_2 _37516_ (.A1(_09541_),
    .A2(_09546_),
    .B1(_09539_),
    .X(_09686_));
 sky130_fd_sc_hd__xnor2_2 _37517_ (.A(_09685_),
    .B(_09686_),
    .Y(_09687_));
 sky130_fd_sc_hd__xor2_2 _37518_ (.A(_09676_),
    .B(_09687_),
    .X(_09688_));
 sky130_fd_sc_hd__a2bb2o_2 _37519_ (.A1_N(_05543_),
    .A2_N(_08931_),
    .B1(_04005_),
    .B2(_00567_),
    .X(_09689_));
 sky130_fd_sc_hd__o21ai_2 _37520_ (.A1(_08926_),
    .A2(_08963_),
    .B1(_09689_),
    .Y(_09690_));
 sky130_fd_sc_hd__a31o_2 _37521_ (.A1(_05450_),
    .A2(_06983_),
    .A3(_08763_),
    .B1(_09532_),
    .X(_09691_));
 sky130_fd_sc_hd__xnor2_2 _37522_ (.A(_09690_),
    .B(_09691_),
    .Y(_09692_));
 sky130_fd_sc_hd__xor2_2 _37523_ (.A(_09688_),
    .B(_09692_),
    .X(_09694_));
 sky130_fd_sc_hd__xnor2_2 _37524_ (.A(_09675_),
    .B(_09694_),
    .Y(_09695_));
 sky130_fd_sc_hd__a21oi_2 _37525_ (.A1(_09550_),
    .A2(_09552_),
    .B1(_09548_),
    .Y(_09696_));
 sky130_fd_sc_hd__xnor2_2 _37526_ (.A(_09554_),
    .B(_09696_),
    .Y(_09697_));
 sky130_fd_sc_hd__or2_2 _37527_ (.A(_09695_),
    .B(_09697_),
    .X(_09698_));
 sky130_fd_sc_hd__nand2_2 _37528_ (.A(_09695_),
    .B(_09697_),
    .Y(_09699_));
 sky130_fd_sc_hd__o211a_2 _37529_ (.A1(_09673_),
    .A2(_09674_),
    .B1(_09698_),
    .C1(_09699_),
    .X(_09700_));
 sky130_fd_sc_hd__a211oi_2 _37530_ (.A1(_09698_),
    .A2(_09699_),
    .B1(_09673_),
    .C1(_09674_),
    .Y(_09701_));
 sky130_fd_sc_hd__or3_2 _37531_ (.A(_09560_),
    .B(_09700_),
    .C(_09701_),
    .X(_09702_));
 sky130_fd_sc_hd__o21ai_2 _37532_ (.A1(_09700_),
    .A2(_09701_),
    .B1(_09560_),
    .Y(_09703_));
 sky130_fd_sc_hd__and2b_2 _37533_ (.A_N(_09565_),
    .B(_09564_),
    .X(_09705_));
 sky130_fd_sc_hd__and2_2 _37534_ (.A(_09445_),
    .B(_09566_),
    .X(_09706_));
 sky130_fd_sc_hd__a211o_2 _37535_ (.A1(_09702_),
    .A2(_09703_),
    .B1(_09705_),
    .C1(_09706_),
    .X(_09707_));
 sky130_fd_sc_hd__inv_2 _37536_ (.A(_09707_),
    .Y(_09708_));
 sky130_fd_sc_hd__o211a_2 _37537_ (.A1(_09705_),
    .A2(_09706_),
    .B1(_09702_),
    .C1(_09703_),
    .X(_09709_));
 sky130_fd_sc_hd__nor2_2 _37538_ (.A(_09708_),
    .B(_09709_),
    .Y(_09710_));
 sky130_fd_sc_hd__o21ba_2 _37539_ (.A1(_09572_),
    .A2(_09577_),
    .B1_N(_09570_),
    .X(_09711_));
 sky130_fd_sc_hd__xnor2_2 _37540_ (.A(_09710_),
    .B(_09711_),
    .Y(_09712_));
 sky130_fd_sc_hd__xnor2_2 _37541_ (.A(_09672_),
    .B(_09712_),
    .Y(_09713_));
 sky130_fd_sc_hd__xnor2_2 _37542_ (.A(_00522_),
    .B(_09713_),
    .Y(_09714_));
 sky130_fd_sc_hd__and3_2 _37543_ (.A(_09642_),
    .B(_09623_),
    .C(_09714_),
    .X(_09716_));
 sky130_fd_sc_hd__nand2_2 _37544_ (.A(_09642_),
    .B(_09623_),
    .Y(_09717_));
 sky130_fd_sc_hd__nor2b_2 _37545_ (.A(_09714_),
    .B_N(_09717_),
    .Y(_09718_));
 sky130_fd_sc_hd__nor2_2 _37546_ (.A(_09716_),
    .B(_09718_),
    .Y(_09719_));
 sky130_fd_sc_hd__xnor2_2 _37547_ (.A(_09641_),
    .B(_09719_),
    .Y(_09720_));
 sky130_fd_sc_hd__xor2_2 _37548_ (.A(_00882_),
    .B(_09720_),
    .X(_09721_));
 sky130_fd_sc_hd__a21oi_2 _37549_ (.A1(_09636_),
    .A2(_09640_),
    .B1(_09634_),
    .Y(_09722_));
 sky130_fd_sc_hd__xnor2_2 _37550_ (.A(_09721_),
    .B(_09722_),
    .Y(oO[91]));
 sky130_fd_sc_hd__o21ai_2 _37551_ (.A1(_09570_),
    .A2(_09709_),
    .B1(_09707_),
    .Y(_09723_));
 sky130_fd_sc_hd__a21oi_2 _37552_ (.A1(_09571_),
    .A2(_09707_),
    .B1(_09709_),
    .Y(_09724_));
 sky130_fd_sc_hd__nor2_2 _37553_ (.A(_09554_),
    .B(_09696_),
    .Y(_09726_));
 sky130_fd_sc_hd__nand2_2 _37554_ (.A(_09688_),
    .B(_09692_),
    .Y(_09727_));
 sky130_fd_sc_hd__a2bb2o_2 _37555_ (.A1_N(_06023_),
    .A2_N(_08931_),
    .B1(_04005_),
    .B2(_08613_),
    .X(_09728_));
 sky130_fd_sc_hd__o21a_2 _37556_ (.A1(_08926_),
    .A2(_09267_),
    .B1(_09728_),
    .X(_09729_));
 sky130_fd_sc_hd__nor2_2 _37557_ (.A(_08926_),
    .B(_08963_),
    .Y(_09730_));
 sky130_fd_sc_hd__o21ai_2 _37558_ (.A1(_09730_),
    .A2(_09691_),
    .B1(_09689_),
    .Y(_09731_));
 sky130_fd_sc_hd__xnor2_2 _37559_ (.A(_09729_),
    .B(_09731_),
    .Y(_09732_));
 sky130_fd_sc_hd__a21o_2 _37560_ (.A1(_09680_),
    .A2(_09681_),
    .B1(_09678_),
    .X(_09733_));
 sky130_fd_sc_hd__nor2_2 _37561_ (.A(_04782_),
    .B(_08394_),
    .Y(_09734_));
 sky130_fd_sc_hd__xor2_2 _37562_ (.A(_09677_),
    .B(_09734_),
    .X(_09735_));
 sky130_fd_sc_hd__nor2_2 _37563_ (.A(_08582_),
    .B(_07983_),
    .Y(_09737_));
 sky130_fd_sc_hd__xnor2_2 _37564_ (.A(_09735_),
    .B(_09737_),
    .Y(_09738_));
 sky130_fd_sc_hd__o211a_2 _37565_ (.A1(_09264_),
    .A2(_09683_),
    .B1(_08613_),
    .C1(_06783_),
    .X(_09739_));
 sky130_fd_sc_hd__xnor2_2 _37566_ (.A(_09738_),
    .B(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__xor2_2 _37567_ (.A(_09733_),
    .B(_09740_),
    .X(_09741_));
 sky130_fd_sc_hd__xnor2_2 _37568_ (.A(_09732_),
    .B(_09741_),
    .Y(_09742_));
 sky130_fd_sc_hd__xor2_2 _37569_ (.A(_09727_),
    .B(_09742_),
    .X(_09743_));
 sky130_fd_sc_hd__and2b_2 _37570_ (.A_N(_09685_),
    .B(_09686_),
    .X(_09744_));
 sky130_fd_sc_hd__a21oi_2 _37571_ (.A1(_09676_),
    .A2(_09687_),
    .B1(_09744_),
    .Y(_09745_));
 sky130_fd_sc_hd__xor2_2 _37572_ (.A(_09743_),
    .B(_09745_),
    .X(_09746_));
 sky130_fd_sc_hd__a21boi_2 _37573_ (.A1(_09675_),
    .A2(_09694_),
    .B1_N(_09698_),
    .Y(_09748_));
 sky130_fd_sc_hd__xor2_2 _37574_ (.A(_09746_),
    .B(_09748_),
    .X(_09749_));
 sky130_fd_sc_hd__xnor2_2 _37575_ (.A(_09726_),
    .B(_09749_),
    .Y(_09750_));
 sky130_fd_sc_hd__and2b_2 _37576_ (.A_N(_09700_),
    .B(_09702_),
    .X(_09751_));
 sky130_fd_sc_hd__xnor2_2 _37577_ (.A(_09750_),
    .B(_09751_),
    .Y(_09752_));
 sky130_fd_sc_hd__a311o_2 _37578_ (.A1(_09574_),
    .A2(_09576_),
    .A3(_09723_),
    .B1(_09724_),
    .C1(_09752_),
    .X(_09753_));
 sky130_fd_sc_hd__a31o_2 _37579_ (.A1(_09574_),
    .A2(_09576_),
    .A3(_09723_),
    .B1(_09724_),
    .X(_09754_));
 sky130_fd_sc_hd__nand2_2 _37580_ (.A(_09752_),
    .B(_09754_),
    .Y(_09755_));
 sky130_fd_sc_hd__nand2_2 _37581_ (.A(_09753_),
    .B(_09755_),
    .Y(_09756_));
 sky130_fd_sc_hd__inv_2 _37582_ (.A(_09603_),
    .Y(_09757_));
 sky130_fd_sc_hd__and2b_2 _37583_ (.A_N(_09665_),
    .B(_09664_),
    .X(_09759_));
 sky130_fd_sc_hd__a21oi_2 _37584_ (.A1(_09757_),
    .A2(_09663_),
    .B1(_09759_),
    .Y(_09760_));
 sky130_fd_sc_hd__o21ba_2 _37585_ (.A1(_09653_),
    .A2(_09655_),
    .B1_N(_09658_),
    .X(_09761_));
 sky130_fd_sc_hd__or2b_2 _37586_ (.A(_09662_),
    .B_N(_09661_),
    .X(_09762_));
 sky130_fd_sc_hd__and3_2 _37587_ (.A(iY[61]),
    .B(iX[63]),
    .C(_09582_),
    .X(_09763_));
 sky130_fd_sc_hd__nand2_2 _37588_ (.A(iX[62]),
    .B(iY[62]),
    .Y(_09764_));
 sky130_fd_sc_hd__xor2_2 _37589_ (.A(_09763_),
    .B(_09764_),
    .X(_09765_));
 sky130_fd_sc_hd__a31o_2 _37590_ (.A1(iX[61]),
    .A2(iY[62]),
    .A3(_09651_),
    .B1(_09648_),
    .X(_09766_));
 sky130_fd_sc_hd__xnor2_2 _37591_ (.A(_09765_),
    .B(_09766_),
    .Y(_09767_));
 sky130_fd_sc_hd__nand2_2 _37592_ (.A(iX[61]),
    .B(iY[63]),
    .Y(_09768_));
 sky130_fd_sc_hd__xnor2_2 _37593_ (.A(_09767_),
    .B(_09768_),
    .Y(_09770_));
 sky130_fd_sc_hd__xnor2_2 _37594_ (.A(_09762_),
    .B(_09770_),
    .Y(_09771_));
 sky130_fd_sc_hd__xnor2_2 _37595_ (.A(_09761_),
    .B(_09771_),
    .Y(_09772_));
 sky130_fd_sc_hd__and2b_2 _37596_ (.A_N(_09760_),
    .B(_09772_),
    .X(_09773_));
 sky130_fd_sc_hd__and2b_2 _37597_ (.A_N(_09772_),
    .B(_09760_),
    .X(_09774_));
 sky130_fd_sc_hd__nor2_2 _37598_ (.A(_09773_),
    .B(_09774_),
    .Y(_09775_));
 sky130_fd_sc_hd__o31a_2 _37599_ (.A1(_09613_),
    .A2(_09619_),
    .A3(_09667_),
    .B1(_09668_),
    .X(_09776_));
 sky130_fd_sc_hd__xor2_2 _37600_ (.A(_09775_),
    .B(_09776_),
    .X(_09777_));
 sky130_fd_sc_hd__xor2_2 _37601_ (.A(_09756_),
    .B(_09777_),
    .X(_09778_));
 sky130_fd_sc_hd__or2b_2 _37602_ (.A(_00924_),
    .B_N(_09778_),
    .X(_09779_));
 sky130_fd_sc_hd__or2b_2 _37603_ (.A(_09778_),
    .B_N(_00924_),
    .X(_09781_));
 sky130_fd_sc_hd__nand2_2 _37604_ (.A(_09779_),
    .B(_09781_),
    .Y(_09782_));
 sky130_fd_sc_hd__and2b_2 _37605_ (.A_N(_09672_),
    .B(_09712_),
    .X(_09783_));
 sky130_fd_sc_hd__a21oi_2 _37606_ (.A1(_00522_),
    .A2(_09713_),
    .B1(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__or2_2 _37607_ (.A(_09782_),
    .B(_09784_),
    .X(_09785_));
 sky130_fd_sc_hd__nand2_2 _37608_ (.A(_09782_),
    .B(_09784_),
    .Y(_09786_));
 sky130_fd_sc_hd__and2_4 _37609_ (.A(_09785_),
    .B(_09786_),
    .X(_09787_));
 sky130_fd_sc_hd__and3_4 _37610_ (.A(_09384_),
    .B(_09391_),
    .C(_09517_),
    .X(_09788_));
 sky130_fd_sc_hd__nand2b_2 _37611_ (.A_N(_09717_),
    .B(_09714_),
    .Y(_09789_));
 sky130_fd_sc_hd__a21o_2 _37612_ (.A1(_09626_),
    .A2(_09789_),
    .B1(_09718_),
    .X(_09790_));
 sky130_fd_sc_hd__or2_4 _37613_ (.A(_09631_),
    .B(_09790_),
    .X(_09792_));
 sky130_fd_sc_hd__a21o_2 _37614_ (.A1(_09629_),
    .A2(_09719_),
    .B1(_09790_),
    .X(_09793_));
 sky130_fd_sc_hd__o21ai_2 _37615_ (.A1(_09788_),
    .A2(_09792_),
    .B1(_09793_),
    .Y(_09794_));
 sky130_fd_sc_hd__xnor2_2 _37616_ (.A(_09787_),
    .B(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__xor2_2 _37617_ (.A(_01299_),
    .B(_09795_),
    .X(_09796_));
 sky130_fd_sc_hd__nor2_2 _37618_ (.A(_00882_),
    .B(_09720_),
    .Y(_09797_));
 sky130_fd_sc_hd__nand2_2 _37619_ (.A(_00882_),
    .B(_09720_),
    .Y(_09798_));
 sky130_fd_sc_hd__o21a_2 _37620_ (.A1(_09634_),
    .A2(_09797_),
    .B1(_09798_),
    .X(_09799_));
 sky130_fd_sc_hd__a31o_2 _37621_ (.A1(_09636_),
    .A2(_09640_),
    .A3(_09721_),
    .B1(_09799_),
    .X(_09800_));
 sky130_fd_sc_hd__xor2_2 _37622_ (.A(_09796_),
    .B(_09800_),
    .X(oO[92]));
 sky130_fd_sc_hd__o211a_2 _37623_ (.A1(_09788_),
    .A2(_09792_),
    .B1(_09793_),
    .C1(_09787_),
    .X(_09802_));
 sky130_fd_sc_hd__or2_2 _37624_ (.A(_09750_),
    .B(_09751_),
    .X(_09803_));
 sky130_fd_sc_hd__nor2_2 _37625_ (.A(_09746_),
    .B(_09748_),
    .Y(_09804_));
 sky130_fd_sc_hd__and2_2 _37626_ (.A(_09726_),
    .B(_09749_),
    .X(_09805_));
 sky130_fd_sc_hd__nand2_2 _37627_ (.A(_09732_),
    .B(_09741_),
    .Y(_09806_));
 sky130_fd_sc_hd__a22oi_2 _37628_ (.A1(_09677_),
    .A2(_09734_),
    .B1(_09735_),
    .B2(_09737_),
    .Y(_09807_));
 sky130_fd_sc_hd__or2_2 _37629_ (.A(_08795_),
    .B(_08394_),
    .X(_09808_));
 sky130_fd_sc_hd__nor2_2 _37630_ (.A(_08571_),
    .B(_07983_),
    .Y(_09809_));
 sky130_fd_sc_hd__xnor2_2 _37631_ (.A(_09808_),
    .B(_09809_),
    .Y(_09810_));
 sky130_fd_sc_hd__or2b_2 _37632_ (.A(_09807_),
    .B_N(_09810_),
    .X(_09811_));
 sky130_fd_sc_hd__or2b_2 _37633_ (.A(_09810_),
    .B_N(_09807_),
    .X(_09813_));
 sky130_fd_sc_hd__nand2_2 _37634_ (.A(_09811_),
    .B(_09813_),
    .Y(_09814_));
 sky130_fd_sc_hd__o211a_2 _37635_ (.A1(_09730_),
    .A2(_09691_),
    .B1(_09729_),
    .C1(_09689_),
    .X(_09815_));
 sky130_fd_sc_hd__a31o_2 _37636_ (.A1(_08613_),
    .A2(_07472_),
    .A3(_08763_),
    .B1(_09815_),
    .X(_09816_));
 sky130_fd_sc_hd__o22a_2 _37637_ (.A1(_08582_),
    .A2(_08931_),
    .B1(_08164_),
    .B2(_04782_),
    .X(_09817_));
 sky130_fd_sc_hd__a31o_2 _37638_ (.A1(_07007_),
    .A2(_06154_),
    .A3(_08763_),
    .B1(_09817_),
    .X(_09818_));
 sky130_fd_sc_hd__xor2_2 _37639_ (.A(_09816_),
    .B(_09818_),
    .X(_09819_));
 sky130_fd_sc_hd__xnor2_2 _37640_ (.A(_09814_),
    .B(_09819_),
    .Y(_09820_));
 sky130_fd_sc_hd__xnor2_2 _37641_ (.A(_09806_),
    .B(_09820_),
    .Y(_09821_));
 sky130_fd_sc_hd__or2b_2 _37642_ (.A(_09738_),
    .B_N(_09739_),
    .X(_09822_));
 sky130_fd_sc_hd__a21bo_2 _37643_ (.A1(_09733_),
    .A2(_09740_),
    .B1_N(_09822_),
    .X(_09824_));
 sky130_fd_sc_hd__xnor2_2 _37644_ (.A(_09821_),
    .B(_09824_),
    .Y(_09825_));
 sky130_fd_sc_hd__or2b_2 _37645_ (.A(_09745_),
    .B_N(_09743_),
    .X(_09826_));
 sky130_fd_sc_hd__o21a_2 _37646_ (.A1(_09727_),
    .A2(_09742_),
    .B1(_09826_),
    .X(_09827_));
 sky130_fd_sc_hd__xnor2_2 _37647_ (.A(_09825_),
    .B(_09827_),
    .Y(_09828_));
 sky130_fd_sc_hd__o21ai_2 _37648_ (.A1(_09804_),
    .A2(_09805_),
    .B1(_09828_),
    .Y(_09829_));
 sky130_fd_sc_hd__or3_2 _37649_ (.A(_09804_),
    .B(_09805_),
    .C(_09828_),
    .X(_09830_));
 sky130_fd_sc_hd__nand2_2 _37650_ (.A(_09829_),
    .B(_09830_),
    .Y(_09831_));
 sky130_fd_sc_hd__and3_2 _37651_ (.A(_09803_),
    .B(_09753_),
    .C(_09831_),
    .X(_09832_));
 sky130_fd_sc_hd__a21o_2 _37652_ (.A1(_09803_),
    .A2(_09753_),
    .B1(_09831_),
    .X(_09833_));
 sky130_fd_sc_hd__nor2b_2 _37653_ (.A(_09832_),
    .B_N(_09833_),
    .Y(_09835_));
 sky130_fd_sc_hd__o311a_2 _37654_ (.A1(_09613_),
    .A2(_09619_),
    .A3(_09667_),
    .B1(_09668_),
    .C1(_09775_),
    .X(_09836_));
 sky130_fd_sc_hd__and3_2 _37655_ (.A(_09600_),
    .B(_09661_),
    .C(_09770_),
    .X(_09837_));
 sky130_fd_sc_hd__and2b_2 _37656_ (.A_N(_09761_),
    .B(_09771_),
    .X(_09838_));
 sky130_fd_sc_hd__nand4_2 _37657_ (.A(_09580_),
    .B(_09598_),
    .C(_09661_),
    .D(_09770_),
    .Y(_09839_));
 sky130_fd_sc_hd__a21oi_2 _37658_ (.A1(_09582_),
    .A2(_09764_),
    .B1(_09645_),
    .Y(_09840_));
 sky130_fd_sc_hd__and3_2 _37659_ (.A(iY[62]),
    .B(iX[63]),
    .C(_09840_),
    .X(_09841_));
 sky130_fd_sc_hd__a21oi_2 _37660_ (.A1(iY[62]),
    .A2(iX[63]),
    .B1(_09840_),
    .Y(_09842_));
 sky130_fd_sc_hd__or2_2 _37661_ (.A(_09841_),
    .B(_09842_),
    .X(_09843_));
 sky130_fd_sc_hd__nand2_2 _37662_ (.A(iX[62]),
    .B(iY[63]),
    .Y(_09844_));
 sky130_fd_sc_hd__xnor2_2 _37663_ (.A(_09843_),
    .B(_09844_),
    .Y(_09846_));
 sky130_fd_sc_hd__nand2_2 _37664_ (.A(_09839_),
    .B(_09846_),
    .Y(_09847_));
 sky130_fd_sc_hd__or2_2 _37665_ (.A(_09839_),
    .B(_09846_),
    .X(_09848_));
 sky130_fd_sc_hd__and2_2 _37666_ (.A(_09847_),
    .B(_09848_),
    .X(_09849_));
 sky130_fd_sc_hd__and2b_2 _37667_ (.A_N(_09765_),
    .B(_09766_),
    .X(_09850_));
 sky130_fd_sc_hd__a31oi_2 _37668_ (.A1(iX[61]),
    .A2(iY[63]),
    .A3(_09767_),
    .B1(_09850_),
    .Y(_09851_));
 sky130_fd_sc_hd__xnor2_2 _37669_ (.A(_09849_),
    .B(_09851_),
    .Y(_09852_));
 sky130_fd_sc_hd__o21a_2 _37670_ (.A1(_09837_),
    .A2(_09838_),
    .B1(_09852_),
    .X(_09853_));
 sky130_fd_sc_hd__nor3_2 _37671_ (.A(_09837_),
    .B(_09838_),
    .C(_09852_),
    .Y(_09854_));
 sky130_fd_sc_hd__nor2_2 _37672_ (.A(_09853_),
    .B(_09854_),
    .Y(_09855_));
 sky130_fd_sc_hd__nor3_2 _37673_ (.A(_09773_),
    .B(_09836_),
    .C(_09855_),
    .Y(_09857_));
 sky130_fd_sc_hd__o21a_2 _37674_ (.A1(_09773_),
    .A2(_09836_),
    .B1(_09855_),
    .X(_09858_));
 sky130_fd_sc_hd__or2_2 _37675_ (.A(_09857_),
    .B(_09858_),
    .X(_09859_));
 sky130_fd_sc_hd__buf_6 _37676_ (.A(_09859_),
    .X(_09860_));
 sky130_fd_sc_hd__xor2_2 _37677_ (.A(_09835_),
    .B(_09860_),
    .X(_09861_));
 sky130_fd_sc_hd__xnor2_2 _37678_ (.A(_01334_),
    .B(_09861_),
    .Y(_09862_));
 sky130_fd_sc_hd__o21ai_2 _37679_ (.A1(_09756_),
    .A2(_09777_),
    .B1(_09779_),
    .Y(_09863_));
 sky130_fd_sc_hd__xnor2_2 _37680_ (.A(_09862_),
    .B(_09863_),
    .Y(_09864_));
 sky130_fd_sc_hd__inv_2 _37681_ (.A(_09864_),
    .Y(_09865_));
 sky130_fd_sc_hd__nand2_2 _37682_ (.A(_09785_),
    .B(_09865_),
    .Y(_09866_));
 sky130_fd_sc_hd__and2b_2 _37683_ (.A_N(_09785_),
    .B(_09864_),
    .X(_09868_));
 sky130_fd_sc_hd__inv_2 _37684_ (.A(_09868_),
    .Y(_09869_));
 sky130_fd_sc_hd__o2111ai_4 _37685_ (.A1(_09788_),
    .A2(_09792_),
    .B1(_09793_),
    .C1(_09864_),
    .D1(_09787_),
    .Y(_09870_));
 sky130_fd_sc_hd__o211a_2 _37686_ (.A1(_09802_),
    .A2(_09866_),
    .B1(_09869_),
    .C1(_09870_),
    .X(_09871_));
 sky130_fd_sc_hd__xor2_2 _37687_ (.A(_01506_),
    .B(_09871_),
    .X(_09872_));
 sky130_fd_sc_hd__and2_2 _37688_ (.A(_01299_),
    .B(_09795_),
    .X(_09873_));
 sky130_fd_sc_hd__a21oi_2 _37689_ (.A1(_09796_),
    .A2(_09800_),
    .B1(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__xnor2_2 _37690_ (.A(_09872_),
    .B(_09874_),
    .Y(oO[93]));
 sky130_fd_sc_hd__and2_2 _37691_ (.A(_09796_),
    .B(_09872_),
    .X(_09875_));
 sky130_fd_sc_hd__o21a_2 _37692_ (.A1(_01506_),
    .A2(_09871_),
    .B1(_09873_),
    .X(_09876_));
 sky130_fd_sc_hd__a21o_2 _37693_ (.A1(_01506_),
    .A2(_09871_),
    .B1(_09876_),
    .X(_09878_));
 sky130_fd_sc_hd__a21oi_2 _37694_ (.A1(_09800_),
    .A2(_09875_),
    .B1(_09878_),
    .Y(_09879_));
 sky130_fd_sc_hd__and2b_2 _37695_ (.A_N(_09862_),
    .B(_09863_),
    .X(_09880_));
 sky130_fd_sc_hd__nor2_2 _37696_ (.A(_09880_),
    .B(_09868_),
    .Y(_09881_));
 sky130_fd_sc_hd__and2b_2 _37697_ (.A_N(_09827_),
    .B(_09825_),
    .X(_09882_));
 sky130_fd_sc_hd__and2b_2 _37698_ (.A_N(_09821_),
    .B(_09824_),
    .X(_09883_));
 sky130_fd_sc_hd__o21ba_2 _37699_ (.A1(_09806_),
    .A2(_09820_),
    .B1_N(_09883_),
    .X(_09884_));
 sky130_fd_sc_hd__or2_2 _37700_ (.A(_09814_),
    .B(_09819_),
    .X(_09885_));
 sky130_fd_sc_hd__o22a_2 _37701_ (.A1(_08571_),
    .A2(_08931_),
    .B1(_08164_),
    .B2(_08795_),
    .X(_09886_));
 sky130_fd_sc_hd__a21o_2 _37702_ (.A1(_08763_),
    .A2(_09677_),
    .B1(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__a31o_2 _37703_ (.A1(_07007_),
    .A2(_06154_),
    .A3(_08763_),
    .B1(_09816_),
    .X(_09889_));
 sky130_fd_sc_hd__or2b_2 _37704_ (.A(_09817_),
    .B_N(_09889_),
    .X(_09890_));
 sky130_fd_sc_hd__xnor2_2 _37705_ (.A(_09887_),
    .B(_09890_),
    .Y(_09891_));
 sky130_fd_sc_hd__or3_2 _37706_ (.A(_07983_),
    .B(_08394_),
    .C(_09677_),
    .X(_09892_));
 sky130_fd_sc_hd__xnor2_2 _37707_ (.A(_09891_),
    .B(_09892_),
    .Y(_09893_));
 sky130_fd_sc_hd__a21o_2 _37708_ (.A1(_09811_),
    .A2(_09885_),
    .B1(_09893_),
    .X(_09894_));
 sky130_fd_sc_hd__nand3_2 _37709_ (.A(_09811_),
    .B(_09885_),
    .C(_09893_),
    .Y(_09895_));
 sky130_fd_sc_hd__and2_2 _37710_ (.A(_09894_),
    .B(_09895_),
    .X(_09896_));
 sky130_fd_sc_hd__xnor2_2 _37711_ (.A(_09884_),
    .B(_09896_),
    .Y(_09897_));
 sky130_fd_sc_hd__xnor2_2 _37712_ (.A(_09882_),
    .B(_09897_),
    .Y(_09898_));
 sky130_fd_sc_hd__a21o_2 _37713_ (.A1(_09829_),
    .A2(_09833_),
    .B1(_09898_),
    .X(_09900_));
 sky130_fd_sc_hd__nand3_2 _37714_ (.A(_09829_),
    .B(_09833_),
    .C(_09898_),
    .Y(_09901_));
 sky130_fd_sc_hd__nand2_2 _37715_ (.A(_09900_),
    .B(_09901_),
    .Y(_09902_));
 sky130_fd_sc_hd__nor2_2 _37716_ (.A(_09853_),
    .B(_09858_),
    .Y(_09903_));
 sky130_fd_sc_hd__or2b_2 _37717_ (.A(_09851_),
    .B_N(_09849_),
    .X(_09904_));
 sky130_fd_sc_hd__nand2_2 _37718_ (.A(iX[63]),
    .B(iY[63]),
    .Y(_09905_));
 sky130_fd_sc_hd__o21ba_2 _37719_ (.A1(_09842_),
    .A2(_09844_),
    .B1_N(_09841_),
    .X(_09906_));
 sky130_fd_sc_hd__xnor2_2 _37720_ (.A(_09905_),
    .B(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__a21o_2 _37721_ (.A1(_09848_),
    .A2(_09904_),
    .B1(_09907_),
    .X(_09908_));
 sky130_fd_sc_hd__nand3_2 _37722_ (.A(_09848_),
    .B(_09904_),
    .C(_09907_),
    .Y(_09909_));
 sky130_fd_sc_hd__nand2_2 _37723_ (.A(_09908_),
    .B(_09909_),
    .Y(_09911_));
 sky130_fd_sc_hd__xnor2_2 _37724_ (.A(_09903_),
    .B(_09911_),
    .Y(_09912_));
 sky130_fd_sc_hd__xnor2_2 _37725_ (.A(_09902_),
    .B(_09912_),
    .Y(_09913_));
 sky130_fd_sc_hd__xnor2_2 _37726_ (.A(_01729_),
    .B(_09913_),
    .Y(_09914_));
 sky130_fd_sc_hd__and2_2 _37727_ (.A(_09835_),
    .B(_09860_),
    .X(_09915_));
 sky130_fd_sc_hd__a21oi_2 _37728_ (.A1(_01334_),
    .A2(_09861_),
    .B1(_09915_),
    .Y(_09916_));
 sky130_fd_sc_hd__xor2_2 _37729_ (.A(_09914_),
    .B(_09916_),
    .X(_09917_));
 sky130_fd_sc_hd__inv_2 _37730_ (.A(_09917_),
    .Y(_09918_));
 sky130_fd_sc_hd__a21o_2 _37731_ (.A1(_09870_),
    .A2(_09881_),
    .B1(_09918_),
    .X(_09919_));
 sky130_fd_sc_hd__nand3_2 _37732_ (.A(_09870_),
    .B(_09918_),
    .C(_09881_),
    .Y(_09920_));
 sky130_fd_sc_hd__and2_2 _37733_ (.A(_09919_),
    .B(_09920_),
    .X(_09922_));
 sky130_fd_sc_hd__xor2_2 _37734_ (.A(_02095_),
    .B(_09922_),
    .X(_09923_));
 sky130_fd_sc_hd__and2b_2 _37735_ (.A_N(_09879_),
    .B(_09923_),
    .X(_09924_));
 sky130_fd_sc_hd__and2b_2 _37736_ (.A_N(_09923_),
    .B(_09879_),
    .X(_09925_));
 sky130_fd_sc_hd__nor2_2 _37737_ (.A(_09924_),
    .B(_09925_),
    .Y(oO[94]));
 sky130_fd_sc_hd__or2_2 _37738_ (.A(_09914_),
    .B(_09916_),
    .X(_09926_));
 sky130_fd_sc_hd__a21bo_4 _37739_ (.A1(_09882_),
    .A2(_09897_),
    .B1_N(_09900_),
    .X(_09927_));
 sky130_fd_sc_hd__inv_2 _37740_ (.A(_09894_),
    .Y(_09928_));
 sky130_fd_sc_hd__and2b_2 _37741_ (.A_N(_09884_),
    .B(_09896_),
    .X(_09929_));
 sky130_fd_sc_hd__or3_2 _37742_ (.A(_08571_),
    .B(_07983_),
    .C(_09808_),
    .X(_09930_));
 sky130_fd_sc_hd__or2_2 _37743_ (.A(_09891_),
    .B(_09892_),
    .X(_09932_));
 sky130_fd_sc_hd__a2bb2o_2 _37744_ (.A1_N(_08394_),
    .A2_N(_08931_),
    .B1(_04005_),
    .B2(_04451_),
    .X(_09933_));
 sky130_fd_sc_hd__o31a_2 _37745_ (.A1(_07983_),
    .A2(_08394_),
    .A3(_08926_),
    .B1(_09933_),
    .X(_09934_));
 sky130_fd_sc_hd__a2bb2o_2 _37746_ (.A1_N(_09886_),
    .A2_N(_09890_),
    .B1(_08763_),
    .B2(_09677_),
    .X(_09935_));
 sky130_fd_sc_hd__xnor2_2 _37747_ (.A(_09934_),
    .B(_09935_),
    .Y(_09936_));
 sky130_fd_sc_hd__a21o_2 _37748_ (.A1(_09930_),
    .A2(_09932_),
    .B1(_09936_),
    .X(_09937_));
 sky130_fd_sc_hd__nand3_2 _37749_ (.A(_09930_),
    .B(_09932_),
    .C(_09936_),
    .Y(_09938_));
 sky130_fd_sc_hd__and2_2 _37750_ (.A(_09937_),
    .B(_09938_),
    .X(_09939_));
 sky130_fd_sc_hd__o21ai_2 _37751_ (.A1(_09928_),
    .A2(_09929_),
    .B1(_09939_),
    .Y(_09940_));
 sky130_fd_sc_hd__o31a_2 _37752_ (.A1(_09928_),
    .A2(_09929_),
    .A3(_09939_),
    .B1(_09940_),
    .X(_09941_));
 sky130_fd_sc_hd__xnor2_2 _37753_ (.A(_09927_),
    .B(_09941_),
    .Y(_09943_));
 sky130_fd_sc_hd__o221a_2 _37754_ (.A1(_09905_),
    .A2(_09906_),
    .B1(_09911_),
    .B2(_09903_),
    .C1(_09908_),
    .X(_09944_));
 sky130_fd_sc_hd__xnor2_2 _37755_ (.A(_09943_),
    .B(_09944_),
    .Y(_09945_));
 sky130_fd_sc_hd__xnor2_2 _37756_ (.A(_02506_),
    .B(_09945_),
    .Y(_09946_));
 sky130_fd_sc_hd__and3_2 _37757_ (.A(_09900_),
    .B(_09901_),
    .C(_09912_),
    .X(_09947_));
 sky130_fd_sc_hd__a21oi_2 _37758_ (.A1(_01729_),
    .A2(_09913_),
    .B1(_09947_),
    .Y(_09948_));
 sky130_fd_sc_hd__xor2_2 _37759_ (.A(_09946_),
    .B(_09948_),
    .X(_09949_));
 sky130_fd_sc_hd__nand3_2 _37760_ (.A(_09926_),
    .B(_09919_),
    .C(_09949_),
    .Y(_09950_));
 sky130_fd_sc_hd__a21o_2 _37761_ (.A1(_09926_),
    .A2(_09919_),
    .B1(_09949_),
    .X(_09951_));
 sky130_fd_sc_hd__and3_2 _37762_ (.A(_02294_),
    .B(_09950_),
    .C(_09951_),
    .X(_09952_));
 sky130_fd_sc_hd__a21oi_2 _37763_ (.A1(_09950_),
    .A2(_09951_),
    .B1(_02294_),
    .Y(_09954_));
 sky130_fd_sc_hd__nor2_2 _37764_ (.A(_09952_),
    .B(_09954_),
    .Y(_09955_));
 sky130_fd_sc_hd__and2_2 _37765_ (.A(_02095_),
    .B(_09922_),
    .X(_09956_));
 sky130_fd_sc_hd__nor2_2 _37766_ (.A(_09956_),
    .B(_09924_),
    .Y(_09957_));
 sky130_fd_sc_hd__xnor2_2 _37767_ (.A(_09955_),
    .B(_09957_),
    .Y(oO[95]));
 sky130_fd_sc_hd__nand3_2 _37768_ (.A(_02294_),
    .B(_09950_),
    .C(_09951_),
    .Y(_09958_));
 sky130_fd_sc_hd__and4b_2 _37769_ (.A_N(_09954_),
    .B(_09875_),
    .C(_09923_),
    .D(_09958_),
    .X(_09959_));
 sky130_fd_sc_hd__and2_2 _37770_ (.A(_09636_),
    .B(_09721_),
    .X(_09960_));
 sky130_fd_sc_hd__and3_2 _37771_ (.A(_09395_),
    .B(_09523_),
    .C(_09960_),
    .X(_09961_));
 sky130_fd_sc_hd__and4bb_2 _37772_ (.A_N(_07945_),
    .B_N(_09237_),
    .C(_09959_),
    .D(_09961_),
    .X(_09962_));
 sky130_fd_sc_hd__and3_2 _37773_ (.A(_09240_),
    .B(_09959_),
    .C(_09961_),
    .X(_09964_));
 sky130_fd_sc_hd__and3b_2 _37774_ (.A_N(_09954_),
    .B(_09923_),
    .C(_09958_),
    .X(_09965_));
 sky130_fd_sc_hd__a21o_2 _37775_ (.A1(_09638_),
    .A2(_09960_),
    .B1(_09799_),
    .X(_09966_));
 sky130_fd_sc_hd__a21o_2 _37776_ (.A1(_09956_),
    .A2(_09958_),
    .B1(_09954_),
    .X(_09967_));
 sky130_fd_sc_hd__a221o_2 _37777_ (.A1(_09878_),
    .A2(_09965_),
    .B1(_09959_),
    .B2(_09966_),
    .C1(_09967_),
    .X(_09968_));
 sky130_fd_sc_hd__nand2_2 _37778_ (.A(_09917_),
    .B(_09949_),
    .Y(_09969_));
 sky130_fd_sc_hd__a21o_2 _37779_ (.A1(_09870_),
    .A2(_09881_),
    .B1(_09969_),
    .X(_09970_));
 sky130_fd_sc_hd__o21a_2 _37780_ (.A1(_09946_),
    .A2(_09948_),
    .B1(_09926_),
    .X(_09971_));
 sky130_fd_sc_hd__a21o_4 _37781_ (.A1(_09946_),
    .A2(_09948_),
    .B1(_09971_),
    .X(_09972_));
 sky130_fd_sc_hd__and2_2 _37782_ (.A(_09929_),
    .B(_09939_),
    .X(_09973_));
 sky130_fd_sc_hd__and2_2 _37783_ (.A(_09927_),
    .B(_09941_),
    .X(_09975_));
 sky130_fd_sc_hd__and3_2 _37784_ (.A(_04451_),
    .B(_06783_),
    .C(_08763_),
    .X(_09976_));
 sky130_fd_sc_hd__o21a_2 _37785_ (.A1(_09976_),
    .A2(_09935_),
    .B1(_09933_),
    .X(_09977_));
 sky130_fd_sc_hd__or2_2 _37786_ (.A(_08926_),
    .B(_09977_),
    .X(_09978_));
 sky130_fd_sc_hd__nand2_2 _37787_ (.A(_09937_),
    .B(_09978_),
    .Y(_09979_));
 sky130_fd_sc_hd__nand2_2 _37788_ (.A(_09928_),
    .B(_09939_),
    .Y(_09980_));
 sky130_fd_sc_hd__mux2_2 _37789_ (.A0(_09978_),
    .A1(_09979_),
    .S(_09980_),
    .X(_09981_));
 sky130_fd_sc_hd__o21ai_2 _37790_ (.A1(_09973_),
    .A2(_09975_),
    .B1(_09981_),
    .Y(_09982_));
 sky130_fd_sc_hd__or3_2 _37791_ (.A(_09973_),
    .B(_09975_),
    .C(_09981_),
    .X(_09983_));
 sky130_fd_sc_hd__nand2_2 _37792_ (.A(_09982_),
    .B(_09983_),
    .Y(_09984_));
 sky130_fd_sc_hd__nand2b_2 _37793_ (.A_N(_09943_),
    .B(_09944_),
    .Y(_09986_));
 sky130_fd_sc_hd__a21boi_2 _37794_ (.A1(_02506_),
    .A2(_09945_),
    .B1_N(_09986_),
    .Y(_09987_));
 sky130_fd_sc_hd__or2_4 _37795_ (.A(_09984_),
    .B(_09987_),
    .X(_09988_));
 sky130_fd_sc_hd__nand2_2 _37796_ (.A(_09984_),
    .B(_09987_),
    .Y(_09989_));
 sky130_fd_sc_hd__nand2_2 _37797_ (.A(_09988_),
    .B(_09989_),
    .Y(_09990_));
 sky130_fd_sc_hd__a21oi_2 _37798_ (.A1(_09970_),
    .A2(_09972_),
    .B1(_09990_),
    .Y(_09991_));
 sky130_fd_sc_hd__and3_2 _37799_ (.A(_09990_),
    .B(_09970_),
    .C(_09972_),
    .X(_09992_));
 sky130_fd_sc_hd__nor2_2 _37800_ (.A(_09991_),
    .B(_09992_),
    .Y(_09993_));
 sky130_fd_sc_hd__xor2_2 _37801_ (.A(_02888_),
    .B(_09993_),
    .X(_09994_));
 sky130_fd_sc_hd__o31ai_4 _37802_ (.A1(_09962_),
    .A2(_09964_),
    .A3(_09968_),
    .B1(_09994_),
    .Y(_09995_));
 sky130_fd_sc_hd__or4_2 _37803_ (.A(_09994_),
    .B(_09962_),
    .C(_09964_),
    .D(_09968_),
    .X(_09997_));
 sky130_fd_sc_hd__and2_2 _37804_ (.A(_09995_),
    .B(_09997_),
    .X(_09998_));
 sky130_fd_sc_hd__buf_1 _37805_ (.A(_09998_),
    .X(oO[96]));
 sky130_fd_sc_hd__a21o_4 _37806_ (.A1(_09970_),
    .A2(_09972_),
    .B1(_09990_),
    .X(_09999_));
 sky130_fd_sc_hd__o21ba_2 _37807_ (.A1(_08926_),
    .A2(_09980_),
    .B1_N(_09977_),
    .X(_10000_));
 sky130_fd_sc_hd__mux2_2 _37808_ (.A0(_09977_),
    .A1(_10000_),
    .S(_09982_),
    .X(_10001_));
 sky130_fd_sc_hd__nand3_4 _37809_ (.A(_09988_),
    .B(_09999_),
    .C(_10001_),
    .Y(_10002_));
 sky130_fd_sc_hd__a21o_2 _37810_ (.A1(_09988_),
    .A2(_09999_),
    .B1(_10001_),
    .X(_10003_));
 sky130_fd_sc_hd__and3b_2 _37811_ (.A_N(_03285_),
    .B(_10002_),
    .C(_10003_),
    .X(_10004_));
 sky130_fd_sc_hd__a21bo_2 _37812_ (.A1(_10002_),
    .A2(_10003_),
    .B1_N(_03285_),
    .X(_10005_));
 sky130_fd_sc_hd__or2b_4 _37813_ (.A(_10004_),
    .B_N(_10005_),
    .X(_10007_));
 sky130_fd_sc_hd__nand2_2 _37814_ (.A(_02888_),
    .B(_09993_),
    .Y(_10008_));
 sky130_fd_sc_hd__nand2_2 _37815_ (.A(_10008_),
    .B(_09995_),
    .Y(_10009_));
 sky130_fd_sc_hd__xnor2_2 _37816_ (.A(_10007_),
    .B(_10009_),
    .Y(oO[97]));
 sky130_fd_sc_hd__and3_4 _37817_ (.A(_09988_),
    .B(_09999_),
    .C(_10001_),
    .X(_10010_));
 sky130_fd_sc_hd__buf_8 _37818_ (.A(_10010_),
    .X(_10011_));
 sky130_fd_sc_hd__xnor2_2 _37819_ (.A(_03693_),
    .B(_10011_),
    .Y(_10012_));
 sky130_fd_sc_hd__a31o_2 _37820_ (.A1(_10008_),
    .A2(_09995_),
    .A3(_10005_),
    .B1(_10004_),
    .X(_10013_));
 sky130_fd_sc_hd__or2_2 _37821_ (.A(_10012_),
    .B(_10013_),
    .X(_10014_));
 sky130_fd_sc_hd__nand2_2 _37822_ (.A(_10012_),
    .B(_10013_),
    .Y(_10015_));
 sky130_fd_sc_hd__and2_2 _37823_ (.A(_10014_),
    .B(_10015_),
    .X(_10017_));
 sky130_fd_sc_hd__buf_1 _37824_ (.A(_10017_),
    .X(oO[98]));
 sky130_fd_sc_hd__xnor2_2 _37825_ (.A(_03869_),
    .B(_10002_),
    .Y(_10018_));
 sky130_fd_sc_hd__buf_8 _37826_ (.A(_10002_),
    .X(_10019_));
 sky130_fd_sc_hd__buf_6 _37827_ (.A(_10019_),
    .X(_10020_));
 sky130_fd_sc_hd__o21ai_2 _37828_ (.A1(_03672_),
    .A2(_10020_),
    .B1(_10014_),
    .Y(_10021_));
 sky130_fd_sc_hd__xnor2_2 _37829_ (.A(_10018_),
    .B(_10021_),
    .Y(oO[99]));
 sky130_fd_sc_hd__inv_2 _37830_ (.A(_04406_),
    .Y(_10022_));
 sky130_fd_sc_hd__buf_12 _37831_ (.A(_10011_),
    .X(_10023_));
 sky130_fd_sc_hd__xnor2_4 _37832_ (.A(_10022_),
    .B(_10023_),
    .Y(_10024_));
 sky130_fd_sc_hd__or2_4 _37833_ (.A(_10012_),
    .B(_10018_),
    .X(_10026_));
 sky130_fd_sc_hd__a2111o_2 _37834_ (.A1(_10008_),
    .A2(_10005_),
    .B1(_10012_),
    .C1(_10018_),
    .D1(_10004_),
    .X(_10027_));
 sky130_fd_sc_hd__a21o_2 _37835_ (.A1(_03672_),
    .A2(_03869_),
    .B1(_10019_),
    .X(_10028_));
 sky130_fd_sc_hd__and2_2 _37836_ (.A(_10027_),
    .B(_10028_),
    .X(_10029_));
 sky130_fd_sc_hd__o31a_2 _37837_ (.A1(_09995_),
    .A2(_10007_),
    .A3(_10026_),
    .B1(_10029_),
    .X(_10030_));
 sky130_fd_sc_hd__xnor2_2 _37838_ (.A(_10024_),
    .B(_10030_),
    .Y(oO[100]));
 sky130_fd_sc_hd__xnor2_2 _37839_ (.A(_04751_),
    .B(_10011_),
    .Y(_10031_));
 sky130_fd_sc_hd__nor2_2 _37840_ (.A(_10022_),
    .B(_10020_),
    .Y(_10032_));
 sky130_fd_sc_hd__and2b_2 _37841_ (.A_N(_10030_),
    .B(_10024_),
    .X(_10033_));
 sky130_fd_sc_hd__nor2_2 _37842_ (.A(_10032_),
    .B(_10033_),
    .Y(_10034_));
 sky130_fd_sc_hd__xnor2_2 _37843_ (.A(_10031_),
    .B(_10034_),
    .Y(oO[101]));
 sky130_fd_sc_hd__xnor2_2 _37844_ (.A(_05091_),
    .B(_10011_),
    .Y(_10036_));
 sky130_fd_sc_hd__nor2_2 _37845_ (.A(_04751_),
    .B(_10020_),
    .Y(_10037_));
 sky130_fd_sc_hd__nand2_2 _37846_ (.A(_04751_),
    .B(_10020_),
    .Y(_10038_));
 sky130_fd_sc_hd__o31a_2 _37847_ (.A1(_10032_),
    .A2(_10033_),
    .A3(_10037_),
    .B1(_10038_),
    .X(_10039_));
 sky130_fd_sc_hd__xor2_2 _37848_ (.A(_10036_),
    .B(_10039_),
    .X(oO[102]));
 sky130_fd_sc_hd__xnor2_2 _37849_ (.A(_05407_),
    .B(_10011_),
    .Y(_10040_));
 sky130_fd_sc_hd__nor2_2 _37850_ (.A(_05091_),
    .B(_10020_),
    .Y(_10041_));
 sky130_fd_sc_hd__a21o_2 _37851_ (.A1(_10036_),
    .A2(_10039_),
    .B1(_10041_),
    .X(_10042_));
 sky130_fd_sc_hd__xor2_2 _37852_ (.A(_10040_),
    .B(_10042_),
    .X(oO[103]));
 sky130_fd_sc_hd__xnor2_2 _37853_ (.A(_05751_),
    .B(_10023_),
    .Y(_10044_));
 sky130_fd_sc_hd__nand4_2 _37854_ (.A(_10024_),
    .B(_10031_),
    .C(_10036_),
    .D(_10040_),
    .Y(_10045_));
 sky130_fd_sc_hd__or3_4 _37855_ (.A(_10007_),
    .B(_10026_),
    .C(_10045_),
    .X(_10046_));
 sky130_fd_sc_hd__a41o_2 _37856_ (.A1(_10022_),
    .A2(_04751_),
    .A3(_05091_),
    .A4(_05407_),
    .B1(_10019_),
    .X(_10047_));
 sky130_fd_sc_hd__a21o_2 _37857_ (.A1(_10027_),
    .A2(_10028_),
    .B1(_10045_),
    .X(_10048_));
 sky130_fd_sc_hd__o211a_2 _37858_ (.A1(_09995_),
    .A2(_10046_),
    .B1(_10047_),
    .C1(_10048_),
    .X(_10049_));
 sky130_fd_sc_hd__nor2_2 _37859_ (.A(_10044_),
    .B(_10049_),
    .Y(_10050_));
 sky130_fd_sc_hd__and2_2 _37860_ (.A(_10044_),
    .B(_10049_),
    .X(_10051_));
 sky130_fd_sc_hd__nor2_2 _37861_ (.A(_10050_),
    .B(_10051_),
    .Y(oO[104]));
 sky130_fd_sc_hd__xnor2_2 _37862_ (.A(_05912_),
    .B(_10002_),
    .Y(_10052_));
 sky130_fd_sc_hd__buf_8 _37863_ (.A(_10023_),
    .X(_10054_));
 sky130_fd_sc_hd__buf_8 _37864_ (.A(_10054_),
    .X(_10055_));
 sky130_fd_sc_hd__buf_8 _37865_ (.A(_10055_),
    .X(_10056_));
 sky130_fd_sc_hd__a21oi_2 _37866_ (.A1(_05751_),
    .A2(_10056_),
    .B1(_10050_),
    .Y(_10057_));
 sky130_fd_sc_hd__xnor2_2 _37867_ (.A(_10052_),
    .B(_10057_),
    .Y(oO[105]));
 sky130_fd_sc_hd__xnor2_2 _37868_ (.A(_06357_),
    .B(_10002_),
    .Y(_10058_));
 sky130_fd_sc_hd__o21a_2 _37869_ (.A1(_05751_),
    .A2(_05912_),
    .B1(_10054_),
    .X(_10059_));
 sky130_fd_sc_hd__o22a_2 _37870_ (.A1(_05912_),
    .A2(_10056_),
    .B1(_10050_),
    .B2(_10059_),
    .X(_10060_));
 sky130_fd_sc_hd__xor2_2 _37871_ (.A(_10058_),
    .B(_10060_),
    .X(oO[106]));
 sky130_fd_sc_hd__xnor2_4 _37872_ (.A(_06650_),
    .B(_10023_),
    .Y(_10061_));
 sky130_fd_sc_hd__and2_2 _37873_ (.A(_06357_),
    .B(_10054_),
    .X(_10063_));
 sky130_fd_sc_hd__a21o_2 _37874_ (.A1(_10058_),
    .A2(_10060_),
    .B1(_10063_),
    .X(_10064_));
 sky130_fd_sc_hd__xor2_2 _37875_ (.A(_10061_),
    .B(_10064_),
    .X(oO[107]));
 sky130_fd_sc_hd__and4b_4 _37876_ (.A_N(_10044_),
    .B(_10052_),
    .C(_10058_),
    .D(_10061_),
    .X(_10065_));
 sky130_fd_sc_hd__inv_2 _37877_ (.A(_10065_),
    .Y(_10066_));
 sky130_fd_sc_hd__nor2_2 _37878_ (.A(_06650_),
    .B(_10019_),
    .Y(_10067_));
 sky130_fd_sc_hd__a311oi_2 _37879_ (.A1(_10058_),
    .A2(_10059_),
    .A3(_10061_),
    .B1(_10067_),
    .C1(_10063_),
    .Y(_10068_));
 sky130_fd_sc_hd__o21a_2 _37880_ (.A1(_10049_),
    .A2(_10066_),
    .B1(_10068_),
    .X(_10069_));
 sky130_fd_sc_hd__xnor2_2 _37881_ (.A(_06780_),
    .B(_10019_),
    .Y(_10070_));
 sky130_fd_sc_hd__and2b_2 _37882_ (.A_N(_10069_),
    .B(_10070_),
    .X(_10071_));
 sky130_fd_sc_hd__and2b_2 _37883_ (.A_N(_10070_),
    .B(_10069_),
    .X(_10073_));
 sky130_fd_sc_hd__nor2_2 _37884_ (.A(_10071_),
    .B(_10073_),
    .Y(oO[108]));
 sky130_fd_sc_hd__xnor2_2 _37885_ (.A(_07195_),
    .B(_10019_),
    .Y(_10074_));
 sky130_fd_sc_hd__a21oi_2 _37886_ (.A1(_06780_),
    .A2(_10056_),
    .B1(_10071_),
    .Y(_10075_));
 sky130_fd_sc_hd__xnor2_2 _37887_ (.A(_10074_),
    .B(_10075_),
    .Y(oO[109]));
 sky130_fd_sc_hd__xnor2_2 _37888_ (.A(_07429_),
    .B(_10002_),
    .Y(_10076_));
 sky130_fd_sc_hd__o21a_2 _37889_ (.A1(_06780_),
    .A2(_07195_),
    .B1(_10023_),
    .X(_10077_));
 sky130_fd_sc_hd__o22a_2 _37890_ (.A1(_07195_),
    .A2(_10055_),
    .B1(_10071_),
    .B2(_10077_),
    .X(_10078_));
 sky130_fd_sc_hd__and2_2 _37891_ (.A(_10076_),
    .B(_10078_),
    .X(_10079_));
 sky130_fd_sc_hd__nor2_2 _37892_ (.A(_10076_),
    .B(_10078_),
    .Y(_10080_));
 sky130_fd_sc_hd__nor2_2 _37893_ (.A(_10079_),
    .B(_10080_),
    .Y(oO[110]));
 sky130_fd_sc_hd__xnor2_2 _37894_ (.A(_07676_),
    .B(_10002_),
    .Y(_10082_));
 sky130_fd_sc_hd__and2_2 _37895_ (.A(_07429_),
    .B(_10023_),
    .X(_10083_));
 sky130_fd_sc_hd__nor2_2 _37896_ (.A(_10083_),
    .B(_10079_),
    .Y(_10084_));
 sky130_fd_sc_hd__xnor2_2 _37897_ (.A(_10082_),
    .B(_10084_),
    .Y(oO[111]));
 sky130_fd_sc_hd__xnor2_2 _37898_ (.A(_07911_),
    .B(_10054_),
    .Y(_10085_));
 sky130_fd_sc_hd__and2_2 _37899_ (.A(_10076_),
    .B(_10082_),
    .X(_10086_));
 sky130_fd_sc_hd__nand4_4 _37900_ (.A(_10070_),
    .B(_10065_),
    .C(_10074_),
    .D(_10086_),
    .Y(_10087_));
 sky130_fd_sc_hd__or3_4 _37901_ (.A(_09995_),
    .B(_10046_),
    .C(_10087_),
    .X(_10088_));
 sky130_fd_sc_hd__a21o_2 _37902_ (.A1(_10048_),
    .A2(_10047_),
    .B1(_10087_),
    .X(_10089_));
 sky130_fd_sc_hd__nand3_2 _37903_ (.A(_10070_),
    .B(_10074_),
    .C(_10086_),
    .Y(_10091_));
 sky130_fd_sc_hd__a221o_2 _37904_ (.A1(_07676_),
    .A2(_10054_),
    .B1(_10077_),
    .B2(_10086_),
    .C1(_10083_),
    .X(_10092_));
 sky130_fd_sc_hd__o21ba_2 _37905_ (.A1(_10068_),
    .A2(_10091_),
    .B1_N(_10092_),
    .X(_10093_));
 sky130_fd_sc_hd__and3_4 _37906_ (.A(_10088_),
    .B(_10089_),
    .C(_10093_),
    .X(_10094_));
 sky130_fd_sc_hd__or2_4 _37907_ (.A(_10085_),
    .B(_10094_),
    .X(_10095_));
 sky130_fd_sc_hd__nand2_2 _37908_ (.A(_10085_),
    .B(_10094_),
    .Y(_10096_));
 sky130_fd_sc_hd__and2_2 _37909_ (.A(_10095_),
    .B(_10096_),
    .X(_10097_));
 sky130_fd_sc_hd__buf_1 _37910_ (.A(_10097_),
    .X(oO[112]));
 sky130_fd_sc_hd__xnor2_2 _37911_ (.A(_08146_),
    .B(_10054_),
    .Y(_10098_));
 sky130_fd_sc_hd__a21bo_2 _37912_ (.A1(_07911_),
    .A2(_10056_),
    .B1_N(_10095_),
    .X(_10099_));
 sky130_fd_sc_hd__xnor2_2 _37913_ (.A(_10098_),
    .B(_10099_),
    .Y(oO[113]));
 sky130_fd_sc_hd__xnor2_2 _37914_ (.A(_08343_),
    .B(_10023_),
    .Y(_10101_));
 sky130_fd_sc_hd__o21ai_2 _37915_ (.A1(_07911_),
    .A2(_08146_),
    .B1(_10054_),
    .Y(_10102_));
 sky130_fd_sc_hd__a2bb2o_4 _37916_ (.A1_N(_08146_),
    .A2_N(_10056_),
    .B1(_10095_),
    .B2(_10102_),
    .X(_10103_));
 sky130_fd_sc_hd__xnor2_2 _37917_ (.A(_10101_),
    .B(_10103_),
    .Y(oO[114]));
 sky130_fd_sc_hd__xnor2_2 _37918_ (.A(_08540_),
    .B(_10002_),
    .Y(_10104_));
 sky130_fd_sc_hd__inv_2 _37919_ (.A(_10101_),
    .Y(_10105_));
 sky130_fd_sc_hd__or2_2 _37920_ (.A(_08343_),
    .B(_10019_),
    .X(_10106_));
 sky130_fd_sc_hd__o21ai_2 _37921_ (.A1(_10105_),
    .A2(_10103_),
    .B1(_10106_),
    .Y(_10107_));
 sky130_fd_sc_hd__xor2_2 _37922_ (.A(_10104_),
    .B(_10107_),
    .X(oO[115]));
 sky130_fd_sc_hd__xnor2_2 _37923_ (.A(_08737_),
    .B(_10019_),
    .Y(_10109_));
 sky130_fd_sc_hd__nand2_2 _37924_ (.A(_10101_),
    .B(_10104_),
    .Y(_10110_));
 sky130_fd_sc_hd__or3_2 _37925_ (.A(_10085_),
    .B(_10098_),
    .C(_10110_),
    .X(_10111_));
 sky130_fd_sc_hd__nand2_2 _37926_ (.A(_08540_),
    .B(_10054_),
    .Y(_10112_));
 sky130_fd_sc_hd__o211a_2 _37927_ (.A1(_10102_),
    .A2(_10110_),
    .B1(_10112_),
    .C1(_10106_),
    .X(_10113_));
 sky130_fd_sc_hd__o21a_2 _37928_ (.A1(_10094_),
    .A2(_10111_),
    .B1(_10113_),
    .X(_10114_));
 sky130_fd_sc_hd__xor2_2 _37929_ (.A(_10109_),
    .B(_10114_),
    .X(oO[116]));
 sky130_fd_sc_hd__xnor2_2 _37930_ (.A(_08909_),
    .B(_10023_),
    .Y(_10115_));
 sky130_fd_sc_hd__nor2_2 _37931_ (.A(_10109_),
    .B(_10114_),
    .Y(_10116_));
 sky130_fd_sc_hd__o21bai_2 _37932_ (.A1(_08737_),
    .A2(_10020_),
    .B1_N(_10116_),
    .Y(_10117_));
 sky130_fd_sc_hd__xnor2_2 _37933_ (.A(_10115_),
    .B(_10117_),
    .Y(oO[117]));
 sky130_fd_sc_hd__nand2_2 _37934_ (.A(_09067_),
    .B(_10054_),
    .Y(_10119_));
 sky130_fd_sc_hd__or2_2 _37935_ (.A(_09067_),
    .B(_10023_),
    .X(_10120_));
 sky130_fd_sc_hd__nand2_2 _37936_ (.A(_10119_),
    .B(_10120_),
    .Y(_10121_));
 sky130_fd_sc_hd__a21oi_2 _37937_ (.A1(_08737_),
    .A2(_09070_),
    .B1(_10019_),
    .Y(_10122_));
 sky130_fd_sc_hd__o22a_2 _37938_ (.A1(_08909_),
    .A2(_10056_),
    .B1(_10116_),
    .B2(_10122_),
    .X(_10123_));
 sky130_fd_sc_hd__xnor2_2 _37939_ (.A(_10121_),
    .B(_10123_),
    .Y(oO[118]));
 sky130_fd_sc_hd__nand2_2 _37940_ (.A(_09220_),
    .B(_10054_),
    .Y(_10124_));
 sky130_fd_sc_hd__or2_2 _37941_ (.A(_09220_),
    .B(_10023_),
    .X(_10125_));
 sky130_fd_sc_hd__nand2_2 _37942_ (.A(_10124_),
    .B(_10125_),
    .Y(_10126_));
 sky130_fd_sc_hd__a21bo_2 _37943_ (.A1(_10120_),
    .A2(_10123_),
    .B1_N(_10119_),
    .X(_10128_));
 sky130_fd_sc_hd__xnor2_2 _37944_ (.A(_10126_),
    .B(_10128_),
    .Y(oO[119]));
 sky130_fd_sc_hd__or2_2 _37945_ (.A(_10109_),
    .B(_10115_),
    .X(_10129_));
 sky130_fd_sc_hd__or3_2 _37946_ (.A(_10121_),
    .B(_10126_),
    .C(_10129_),
    .X(_10130_));
 sky130_fd_sc_hd__a311o_2 _37947_ (.A1(_10088_),
    .A2(_10089_),
    .A3(_10093_),
    .B1(_10111_),
    .C1(_10130_),
    .X(_10131_));
 sky130_fd_sc_hd__o21ba_2 _37948_ (.A1(_10113_),
    .A2(_10129_),
    .B1_N(_10122_),
    .X(_10132_));
 sky130_fd_sc_hd__o311a_2 _37949_ (.A1(_10121_),
    .A2(_10126_),
    .A3(_10132_),
    .B1(_10124_),
    .C1(_10119_),
    .X(_10133_));
 sky130_fd_sc_hd__xnor2_2 _37950_ (.A(_09375_),
    .B(_10055_),
    .Y(_10134_));
 sky130_fd_sc_hd__a21oi_4 _37951_ (.A1(_10131_),
    .A2(_10133_),
    .B1(_10134_),
    .Y(_10135_));
 sky130_fd_sc_hd__and3_2 _37952_ (.A(_10134_),
    .B(_10131_),
    .C(_10133_),
    .X(_10136_));
 sky130_fd_sc_hd__nor2_2 _37953_ (.A(_10135_),
    .B(_10136_),
    .Y(oO[120]));
 sky130_fd_sc_hd__xnor2_2 _37954_ (.A(_09507_),
    .B(_10019_),
    .Y(_10138_));
 sky130_fd_sc_hd__a21oi_2 _37955_ (.A1(_09375_),
    .A2(_10056_),
    .B1(_10135_),
    .Y(_10139_));
 sky130_fd_sc_hd__xor2_2 _37956_ (.A(_10138_),
    .B(_10139_),
    .X(oO[121]));
 sky130_fd_sc_hd__and2_2 _37957_ (.A(_09621_),
    .B(_10055_),
    .X(_10140_));
 sky130_fd_sc_hd__nor2_2 _37958_ (.A(_09621_),
    .B(_10055_),
    .Y(_10141_));
 sky130_fd_sc_hd__or2_4 _37959_ (.A(_10140_),
    .B(_10141_),
    .X(_10142_));
 sky130_fd_sc_hd__a21oi_2 _37960_ (.A1(_09513_),
    .A2(_09507_),
    .B1(_10020_),
    .Y(_10143_));
 sky130_fd_sc_hd__o2bb2a_2 _37961_ (.A1_N(_09507_),
    .A2_N(_10020_),
    .B1(_10135_),
    .B2(_10143_),
    .X(_10144_));
 sky130_fd_sc_hd__xnor2_2 _37962_ (.A(_10142_),
    .B(_10144_),
    .Y(oO[122]));
 sky130_fd_sc_hd__xnor2_2 _37963_ (.A(_09672_),
    .B(_10055_),
    .Y(_10146_));
 sky130_fd_sc_hd__inv_2 _37964_ (.A(_10142_),
    .Y(_10147_));
 sky130_fd_sc_hd__a21o_2 _37965_ (.A1(_10147_),
    .A2(_10144_),
    .B1(_10140_),
    .X(_10148_));
 sky130_fd_sc_hd__xnor2_2 _37966_ (.A(_10146_),
    .B(_10148_),
    .Y(oO[123]));
 sky130_fd_sc_hd__nand2_2 _37967_ (.A(_09777_),
    .B(_10055_),
    .Y(_10149_));
 sky130_fd_sc_hd__or2_2 _37968_ (.A(_09777_),
    .B(_10055_),
    .X(_10150_));
 sky130_fd_sc_hd__and2_2 _37969_ (.A(_10149_),
    .B(_10150_),
    .X(_10151_));
 sky130_fd_sc_hd__nor2_2 _37970_ (.A(_10142_),
    .B(_10146_),
    .Y(_10152_));
 sky130_fd_sc_hd__and2b_2 _37971_ (.A_N(_10138_),
    .B(_10152_),
    .X(_10153_));
 sky130_fd_sc_hd__o21a_2 _37972_ (.A1(_09621_),
    .A2(_09672_),
    .B1(_10055_),
    .X(_10154_));
 sky130_fd_sc_hd__a221oi_4 _37973_ (.A1(_10143_),
    .A2(_10152_),
    .B1(_10153_),
    .B2(_10135_),
    .C1(_10154_),
    .Y(_10156_));
 sky130_fd_sc_hd__xnor2_2 _37974_ (.A(_10151_),
    .B(_10156_),
    .Y(oO[124]));
 sky130_fd_sc_hd__xnor2_2 _37975_ (.A(_09860_),
    .B(_10055_),
    .Y(_10157_));
 sky130_fd_sc_hd__nor2_2 _37976_ (.A(_09777_),
    .B(_10056_),
    .Y(_10158_));
 sky130_fd_sc_hd__o21a_2 _37977_ (.A1(_10158_),
    .A2(_10156_),
    .B1(_10149_),
    .X(_10159_));
 sky130_fd_sc_hd__xnor2_4 _37978_ (.A(_10157_),
    .B(_10159_),
    .Y(oO[125]));
 sky130_fd_sc_hd__xnor2_2 _37979_ (.A(_09912_),
    .B(_10056_),
    .Y(_10160_));
 sky130_fd_sc_hd__nand2_2 _37980_ (.A(_10151_),
    .B(_10157_),
    .Y(_10161_));
 sky130_fd_sc_hd__o221ai_4 _37981_ (.A1(_09860_),
    .A2(_10020_),
    .B1(_10156_),
    .B2(_10161_),
    .C1(_10149_),
    .Y(_10162_));
 sky130_fd_sc_hd__xor2_2 _37982_ (.A(_10160_),
    .B(_10162_),
    .X(oO[126]));
 sky130_fd_sc_hd__nor2_2 _37983_ (.A(_09912_),
    .B(_10020_),
    .Y(_10164_));
 sky130_fd_sc_hd__a21oi_2 _37984_ (.A1(_10160_),
    .A2(_10162_),
    .B1(_10164_),
    .Y(_10165_));
 sky130_fd_sc_hd__xnor2_2 _37985_ (.A(_09944_),
    .B(_10056_),
    .Y(_10166_));
 sky130_fd_sc_hd__xnor2_4 _37986_ (.A(_10165_),
    .B(_10166_),
    .Y(oO[127]));
 sky130_fd_sc_hd__xnor2_2 _37987_ (.A(_11370_),
    .B(_11385_),
    .Y(oO[32]));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_Left_443 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_Left_442 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_Left_441 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_Left_440 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_Left_439 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_Left_438 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_Left_437 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_Left_436 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_Left_435 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_Left_434 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Left_433 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Left_432 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Left_431 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Left_430 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Left_429 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Left_428 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Left_427 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Left_426 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Left_425 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Left_424 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Left_423 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Left_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Left_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Left_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Left_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Left_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Left_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Left_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Left_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Left_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Left_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Left_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Left_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Left_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Left_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Left_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Left_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Left_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Left_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Left_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Left_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Left_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Left_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Left_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Left_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Left_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Left_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Left_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_Right_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_Right_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_Right_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_Right_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_Right_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_Right_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_Right_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_Right_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_Right_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_Right_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Right_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Right_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Right_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Right_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Right_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Right_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Right_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Right_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Right_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Right_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Right_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Right_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Right_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Right_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Right_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_980 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1095 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_927 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1067 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1094 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1095 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_1265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1094 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_983 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1313 ();
endmodule
